`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Z7wtcnqzGEl1YB6x0obJMp/QqasJsGXn7Ovi+vN+pcuf0Kq9/fsmmFzgWzo2PqsjSidw1UDyOfwD
NJMcBJ25zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TvSSJnXRDTx95zdF03mcP0Nw12huSfiWyui0LS6ZLFjdeo0Pfhv+n2rJavkC3Rp/ZreaLA0XtnLY
rJhjf6642Dq2FQbT7plurVPc8cCLm4aS4orvOJ+Nzv3aRw8UF5gqSlpLdnFsbBl88Xgpjd6DN6vO
hB6bDI3GujhM1pCgEuA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i9/MXTmWw68UYy7En5jmBz+lfIjUO4OkqvGPJqVxTaE0GIBqKseUmxjxrPZEAVLfZYuLDjtGTFFV
xI8JQcBkrlZaCzf4bp78wrAh7st2VujUi9c4ytSmo5PmsSz2IO3gyOw/lOqaYo2YFpHI3pC1Yzce
4JwoJCk/ZVSUfhO+DVAi3y6r6GvPuHNZspcnpolDnbiRZeUrv9gaizfK5afE8qnqMWS4DaEb1WWO
UUn5hZov4ELjgOMCXCjQdEpsX3C8e01yvjD1mK4VZU2cYi+NmZqxOQQy/eDOu3HY0/5uDHqtLGwD
WtJ4DbYcGblTLikRa+3ucLiJhAbNKS+xw/0TVQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zQb7Yu1jeLbG2rH/QGVJyx9WsuufurwlisJ4N5lJs19vc3mFW/MrorYiDBMz8/ZeNbWD9TmO1N15
a6qUT6qawxKXFY/O7hZKIjsVohny35oYjiJp4algKGmiXY6c1zt3ZUbi1z2OccTHSFNMCGIVq3dN
LkJc7cXJl4LqmQqm8fM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BWFO4UcSG4iRfIccMCi7CSeEXuKFkyVMa9CEeM4t23gWAKDtC8AthCnilNOWseLqMDNOu6AchXv7
NevbxD6l6gEL+jczD0lFztdQ61sDcwyKJJhwVlpkP52gErtKxPBejGg8ab9sUv0wCsNt/uTWexST
QKsCcBqIVIDVHJ0Co0jzjBRe++MWa+LU2y94SbJSv5sVC6V2FsumS7IEwUsBkZAbSoMVtQLqsxsy
wjYp/6QVGrRwn0Z9ogpH292TkKG2w9+RUC94IBRwaKWouN4C02nAXuplG6Y6ARvX9ZdgeYTIcXfD
jD/V3wYBt9PMFHEorbEmIj8ZhE53TeoSYVI7zw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gEOGo1TNktG0WMV70jAzFa1dLrb9izaZuDIzmneayRNzUfoCoWD4OzyomeOWT5R7QSFPZG4Noz4J
Kdkl/VhK5dCyS3Hc9BADzqjmkJBLWiXlzv8f+s6Kz4tgjnduDJ+/lPLhAT8YMyAg8dyf9ZObsylp
JNrUQmdVoxA9erwgasXpvfcCnUtC9SGhkD1EYMQTKJfGBIFWcdu6HmtwVZeMry5J1qFHaNKpFxHS
5on14/dcR+rD12bA8M39SnAVl/UDGnlxm3861bAN2lblrWDD87a4Sh1OHsaKaQfXcvLyb1iz4sgC
sGooooUTWU7Lk87EQwMbun8Mu6QRxVWR99hH1Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5904)
`protect data_block
n2C2vFxAn2YB3grmWtGYzoN/EqAH+5lgSstQ1a7+VcGAhV5QCmtGbhCbZFc/ebWRmDrZWHTPuolG
PAYimtSVS/4GDbMELK0H6jnRvslTWSQpPquikYAZXcXxwZ6DgeOAiowGL8Yb9bNqNS/qamvN0jSa
PYJQJpWh1Avpq5FHsDwE600jfERg7TTpNzUdU7JfCFhieMPL4Pz7AcoEvR9hjp2f7ttt9nbm2QHt
251Qm80h4huwD7ahS/s6kLStfgESnT35MJHS77hDhMK8dw+j6fmqzZp41CaCCEFWTTioOJ94oMlR
JLjC5VK1+7pU8kQsi9RzvdSM1ho3NG3AerYWavmy9aRws5RtaM07FhIyHnkqrJ6Qe8EtA1JoMrWX
INGdqR2nQQpQbQK+NoJzUO9XlYGXjNfd90FyOKxQzpOtr6MTCcXAU3EQC3DpnDIwkdayJCbi/cKA
pBuQ+tVVL2nJnZpJzQa39l5o97Y+4NYPG3nCAPIGu62YxOFelZZs2gzqvv+V/KhIrgqh2BDZ0Qqu
ZvGzEDYJiA4tOy+o+sL80TLqZFSbaAGV+LwC00znxP/d1h+MqQYTmhHTiatb+Cwx4e4yK2u+enOc
Y0WGYi+VWqjD2L1oU6pyiod+10go2OE9MaHxFkFJCxtTvIgdx8kkRdSmnJ+oLn9AMnmq8q4n0SNb
ubQAFhj4sTyGvjp7VPqRKE5pPb+/ne2Z17CgiAkVzpnK5Qk+yjw4DsgTXDZTDn7L9NE+AZbz0V8A
5lEmIheyg1JpR8FUPJQ54dM5lLWpEO402uvxdtqfTdMCRpRKG8PoSJ0Ne43VMtRmEutA1bYXkQAf
i3/mDA5/iNP0R4uWHi1UQOIyEVPtCkRMsSVg6iuPSonb1f/xUSZFAksq28JGl1wJZGma328olYGb
1R51oQ6tWY718Xz1GlrVamaaU0VE9BMQp3CIKr82qZpihBN/NSKEFLEcuSxwPvrXf+JmCU2AGfyd
Hbtkwpjt+IrrxcDPXDjs4n82be7Gbvk0bLvZDaA8PN9SpF9MbRNeZuSj+QLgAPCs8kdW/JTQe9sK
keYb+/dChWG3qxtpZ8+ZOnnRYQOgWtkCOt9jTCNWrzQhq9kKVnhzZx3XmaQ58P4H79X7NJlc6rQj
OTcztPazM2ZcxLSxbKFJGplBrcLsL4ITce3Sb5BD1+/appllMUi+dibnL3VEIh6G+wDxJTpzne42
2pz71iSiO/Ti2SWhy8E2tDPa72PhIizB7iF9DDyfg62/g/KrTImSNbqlh2V+wNmH3Xyggndk1A9f
Ugh3L4OGRd1M102HWbSgha8rufsnSzmvkwmDYaA91QfOY15oUYeVhZi8AQOmjoknYWDhQumZkMI6
pSkoAugTKPJIOtyKQvHuvDKPQ+f4cUE3LukOKrc5j9xKewWTeQEhA+5bcxsRnHhSCjt5K3NSz0TM
Qc6o44Nrbvo/uDPYWUXGf6oRMW9C6OxDsAGGql2J5L9MjnRcB53qmcf9kvq5ruFwi2vWzk2rlkvi
/kz13BOqNXGph6RR/IHzT2HPSEduFFBzjzUspwpjmDLxf87iPtzFvqNl1r5wEuJYBot/H4avL4VO
cg+2F1brU3X3KoOKWxJzhSP+AhVwW6c6qE1rpHdwwmMensijmI6vZCv28tC1rrwOzdXcDVu+xtyo
PJ5ETq8ve3ot9pQggZbJA8aICSCDIvSY+mRGhxiVWC1bEd6emn2CSpSp7yfvM5HpjDXRXvtKJekA
DuV6p2HhnUQLRoyTpz4WUfXGWsqFYXOWwH8QwmFwQCfVJS5Tcc4hTS4BNOItfu73W5N+XNX2X+mh
2qKAwdzf+ZZ3Mti1nSGdpyUqmK138qT1kZ7q3dMrQTvZT39TMKAPs1y59hWpuF2FJE6B7TJJzaM1
M2yWLBoC6pqVS5RTaqTr2w16VxJg3JuyO8xbxu1cmwl1uCUCsRxWCqkUXg/N1xkWUSNYXCklFC3F
xRtK3We8GnWittknC0+62MexClfknV2WUzMWzkTzchXokK2x6CkuJbtPaiSUiwnL1jY4toeRr2kr
Kmge+f7iTqAdYy0hHBMOFNbBn+D7Dv/nQT4GvlchFB8mDZBE93l7EJpL8UETflC0pKxkUpMw5gum
M30+V99NDBH3w5cWBZmTlJiDe5u0xHkwIYMSsDWsiY3Q1sYjZZrmsCUWrL5HSbRvB1zhXNNI3YDF
zgvg4nRWxLB1LUmCzBUA3AQDs1REQOijL1pg7o8iEFfJlm2vKdF25H59OeLP1GMPgzz4pgypU7Di
sF5Griw6SM5tcjTnBHKYFINYLWBrTWtT8wheAzhfwkKrB9ynOYvQ66ylcWj95pZkdU9QeTi4OuTB
IztPDM7RdtSOCoIgI2TKd/4Ao+cA3Gbp/S6OcGe7BAdTE5d9MNdoGYSHCLMASn97xBrAGoDmWCBq
6wVCZNILCDWwvFE4hK0M23cwA1AlNDjFWQSU69qdY6XEqdBQw1Qs2QkdoOUVG4/iRkS297Ka4sJh
hmf5mQwHZF5X8BSNKS5ygx/rEe7hHbKvBNlpecJaK/DD6ug1c+dIMm7mKBo+UalR2fB11XMNXjiV
FVs9RGser+R+Ceeww+16axdm1pnth+hVw+E/nWN3GVi3A/5llSufIPGa3Fg/ySWlZMwRJsoH405y
2v9Dxodgn+SyW4KXTmFqsW+3kJ2dfxzOLZzZ2hjy6N3enpHRNAsPfsZMWaXy/3j2NN73a4EcwnkR
4d/90plSRUy26unBCtlItu2luHDzvWyFn/uyGeU66KKB3VhE7MnmZO4VjtgxOPRjRz1sGTs1/p8F
b7DAdEZz0s6W9zFktx/0ZpLvAQhblQYRuko+1Bvw1jb1fIw27gIoIAad0MPe+Gyj1XZR+EJVrv83
6ueBAttxQK+2263fAmRDmJkjUA1tP5Qrw8xx6ml/C6Hsu4AgKL9flM7+zRWwM11EujiYHJi/QJ+c
2unnb6vFVvQ7O1g3P6AWk2jCrmNibomLvU5B5hbes22xdLeSlmv3HJwPTAHn8lFTvWwXRTJ/dCIp
o/YN3Ryo5OFb6GPza7/wcoFniwpPw+aKPRWbbRuQB6pnSQTQ/UWYFvrKRPEpyzJ1e3BZX51j69lp
Z6HWotW25zYPFDI0c1VbdlE61QzLIu5P51lHq9OvEJ4dVnSKxevHlxT/kowsBDyOjzkLEwqc/4RF
Ov0WRFun61JewsINAaw21xSwax1mLIXBY70yQTyvbOPQQ0HoT/6Qlk8E3yPdhEDs9WFGzYy8qx6u
DjQDCAewpDtSq7ySCV1vyfkAsc6JOQwvxZCdsrCVqT/Wtlhapal1/X9HewPSelhy4lhJ6rc60REa
GfpI7joRXmwvBq8EXtMEb4Asutf/ytD3Xz2RkFKmGAxjH6iajxjR2jkvE12H6kl2E36N8fBQ6f5Z
oBZg47aBpQMKeoY1ZM+47+2556pS0hMYCS1gN8Xj6fvgxQ66m3WbSRXi9zeqAOU2th/Qi+VbF16E
emZSo+lPROeUVF8+Hy+dL0L6BJIi5iw0Aj2SGvjTx4ELBlDf6cu8Dt/NfKPqpY+k1Rl7DYJ/6kAR
AELPhZsRTc+8G2aA4gPYrH7Td2B5uj6hLIuvItvNAjUNH0/kGf1X6Dhl1RZwefnmhAeK3i2SXzy+
DrgiQY+gYYg7nAIE2kVqSyzLn1sEHqD1xdpThetW3kH7eQsrFkqh8zP/PtFniz9OmtMxji7pwsE7
ihN876O2xvtMAKfhEurONxBMaIlc5mtJttJTs9NJ+Y9ct/d3eJciJ4DV7/n1cSWyfjeBYJZ+3Uk8
cJbyjWz1LqtSBFPE4eZ5f0GlHDGU3psPMpdgGGzUSJ/DZ4dyDq8uW1Ymyl5v0C9vkzSYgkweidjX
XWM8QUThIlELLadEjSTDc7oQUbgBaO+7sQQHXjYzU4NWjw4lBQmeNC8KZIXp6WfsV2Eu+ZPPnOvV
39u5veSA84pnW0vpKphcqgkVPJS2lYSCJ377ViraTd7n165C/Y3yTuGMFtJ6g4/7C6DDRSg/iDCa
APjKxZIF16PqaknpP5016HDoZObyl//kiCSBVcQpngtsQoxgLjk23eb7foxIoTUKlxNsEQ5rHJfd
4UjNuTY86ZByClYEReLJbr7uPOOL2ddm7tjE35kEgdYxesLT9ru8Y03YA6T7A3dViq3dSiPT5dNu
c5UQGfFamZc65A6SYH5jGJTdwcu7Iv82mwPccUTDpLz2v5exwQ+E/TnkAOV0tmMFIntrCpbMTIvj
7lvy3l4pwQwVWcOx6rW9YvdJT4t/+1qWMr9WO1NVtt0XQio83nkAuAALZfA0JchRPubYpCDt+iDd
MJBNcttOmym/CiEkRHVYK7IKjZltl0eDPfxYwqrzN3H9yBOtVyFdR9EwiY7eoCOzNfSuw9mn839q
JUIbYxYnSotIhO5DZke+ewAsXKpBprdT+ZYLLwcqk9IXlVwCTVZH5tMHLGWKzPlwKr2fGo/NtO+M
VccaHcGA8QxYhQnTdseqASsp5GIrWDl1tCyMhimFVMjPvnFGHIsmXXw9Z4xL7DFTnFOObVTGxq0g
tvGbSgc3qyi5EHGF4EMRk1dXoRg7xl7zh/AZQZCw3DLuGjKb3orQc9vXD2cyhJcOJJcx2mTxEnz3
jafqntg3vAvhGJkxPZvHODwg776ODautNPxWFKzgnIevWsiqZFw6IY8F9EtynnwoT9i46YCLixgD
zg5+JJkYMxyIobtgnWisu8bqpsr/bRz/mb+BkIqbuDJ+x2eMCi47unmpl9JHGJ05mprIP7YNNShj
0NleTrWee3Wxd8Fn1DBNXdUPCUHd1F6XOylx5RfZNJ0McE/8/gfjTGdx50qV7Ad597zxp+hkV9nO
iJ/uwyCMtOkrIckr0rd97gfoTMNpg4UPfgi81OQlGkqDPZbHKvdND1JmGDrbukBGQocYYE/lFCzl
QYwEGlZPRdr5koWcyM6sIFgfrapi8p7DbgEcsHrTACnaUfBuOBCBOjqq9p9bExsG3kL8BzRHMAqT
+qfGo2e8LHgu4kQr+OD5VcngoiNznP30Wbb6EsCPiDw9+s8Gx8uZVkQOJdMCtU/WNSn4Z94vxirW
VNLsrTElr5GosETdyw0armrGISgp+jJ9b7g+cqOXffAWIUN8qI9iKDTqJ+KeyhxDDp6YVSclYVGb
iFsJmMqtURk03V+Lzpz7wV6xai26wPBkam767f5pSnvhFowd5aX7N/Iohb/etNuNyuXn+zJEWRfL
u8xqY9SWIbV3KlR8B5KOURoVOCUJfh+ZE1bjeRYtLZkzg7Bn5WqSivxIKb+zySaR3npXIrHVdwIO
qQZ3D8N090WXdPEa6BHvpt46X5Ffxsg3GhZpt1YTp7a6DGw8E48JphjxNksHl8NxEcBHN6D32w5+
JBb8/zMNQVzUkMm59/gC5pfrne1QkHkYNjRDFXaeqj0ZHpiDwSW3Fi/OQagP6zPzKjcw8zSvjYOU
bqhbOEXpW54W5M/KABOUACMfMBBXqRUJLTpsYB/3POc62tqEvv1gCaRGjvKhYxs8F4ft97o1yaoH
FD9GX9pOlJZA14gjOJBK9PajTwb2TQ7p6FcXjN+kcIgJwBycm0Z2zFRUCEkZiMTW6OWteetJAJ8f
G5TAg+kKRY9ybtw9Rt5GNzTrYCoUW/2q2SnDpqh3U4lurqKIJvmdZwU+fcHsmE4EMHAhYV77o2rL
0X0CjqrFYKq4KQY5XzBEPUrAv0GkE3W/I39Mj3hjvcxgyyxcTEjLbSazcJvRQQsqFqeQqcby5CKj
yaIYo8XMVTQLZqrhPfAaFySVw2EFW8ZbmdqJrnARSMi22I6aFH/tlW+eegpbsrPr7Ld9qn9CEhgF
RMiyyZmzbK8IiicX4ezB8WD6+FWR6LnsnkGZqwx6N3Dsg3aCWkaEKHgK3/iJO/4kziqAR3eTO9XC
DPNwR6XSgRn6U917tutJ7nkknQvb5MsLtF/bGgotAIELhog00FxP4rES1uNcm06zboM2m0S+dKal
rBCvFs5lU9vKrkD5FSQejA7Nx22bpqrFCC9GWh1hQvzhbT0CwCt5G28mtDwGvvjMFvQ4+w0rRREW
R1OuvCSuXXru3nDYUEn7TZYleUhee4VNNpn1tkcNxA3JImiOn6ld/bYyrDNmCYxwrGMsIFzUyzR+
q3PepwzSAOfZxBkvrZpLA2DjiFnxOWGvSyG6NqJSvk2AOZ+BRxA9xQVQBA2JhARTDrrHMtG9X0ME
BtSYzcf8ZQ3kbE9UPBsdd/39f89d/ImPXPK7yH6YPW7qaJ8xHeYvkOSUWilxEtg5wsXqk3B7c761
gq7JOKDHruG0+IvotyBqBK1NR2XnIBok8Zvy2gpbPDFLGv/Bv/B4yqYhSFXoeGTV2aU9iqgHRPz9
uhp1rNq8EZ5lgy1iGCnxJllQZ7mnLlnP8+RUG2YEtns1jZER4RGCnqUNgByrLe/rwDVKxFDiEuVJ
thgtC1P1npsDgcHnajipBX257GCobh7UAltMIVfAgQIjK1deskX2IbEbmhtFIOdLW2rj7gNCixmJ
rftUJjANSKA1Sq1pxOXPaE5o2Eu9qsxrmGLrB+tO34c6+1EyZLPRXiUmeeo9A/j/4Z8fBfEkFfOR
fGjL48JhJvT6HEiZxJHgfFSy4XDZ+HsXHR5gL7PE/PHQS0AaIjLS7m8t5b3K1CFvXXCZfJguR9Ck
YNilaCkb1SAn7z3jioleMlECPTjVxNpek4upvKLbxfvXl2o6yb7cT734Qu6sJTYCIpaOQxHnnKU5
NZb6egAuzsqr/8nD0NO0k6zAevtr3UQH3AFYNMVQllrCMEZSauWTraixrjhVkIo0LJP6Dr8ha0Dd
yeQZ3BbBHwNYpINoqmwSsJzQkr31z2q3t1rlG2uNpDLMvdQAMyxvZl27otBizCVrm15AjSSckWJc
JPBygKql/i3vkJuU7CUs4fyvUUjcJ3p745y269sWys5hQXVfIBVSE3mDATR0rdIszXcvprO8TyAo
Tqss7b9QklexKCwpdnCfVEDMIWU6cLhAmBfSoUuS4ukfHIKNoCCXapJlS9DM/j9cpuvJe2pJUtVX
7b85fQVhOGcphj24hpRYY05540M3CC6Se/HKQuynq9j2LfQ/wog5VUNY7jUkMVs3jOyhqrryMPlz
wUDDfGr5MwdwlkdaGfYRN88V5UfzudZJSAaYyhD0y437xFC3ydmq7mFeO8feNqw9wPO4xSUXjY1J
pALdozTEqWpRuxwDk6w1iHIKqeb0PwQ/nPHK83ydMXqwxLxRTf2ee9owrfnqXuNLUjNwrqtscwb4
1lx5ssOhrygTDsj0N6cGyDIqEY+dpMKDGc/n8p/JfttUYTuysai4gstFOpqeqD6xGvR51t+sBr62
+YUTgPurZ9WGmU/F/Wu7Y7GNIxIKwnxdGRKrjS1V8g0zulmbQ4fLDPBExEOCPhn9+EwwngJfXEDc
MVuMqXsQtOVjqUsNLr+PQ2tGIhzhUIuOdS3u12h0egff3hTT1L+wAq5D4FUbD8Q9CRKqT5j9RUWK
fGU7kDfFp/EGoe4eI9bOJVtWR8R8l2F+4vle64w3uSLOROUeYoVZoAHUwZ2lesPhmFasp6c/9rku
OJBMTeW0e1wI4lm+xtiBGqpM23j2Shp5vfEAUeC5ZzNsrilrVQ8MMyk07n2WCcUw8NUDccR/Bq9L
uZpskBSb2m3L4XQrUx2sOjWToZ9ZMpN18oCsvSR97bUi3ML/+CPrCNHDM+BJ3iIKaXurAatmMMVI
KbgafnI7qHqnYPV8x2gU1RP9EcUPilzuCIS+gs3S2pBeG2Ru1qTnLxrq3b8R9HAOkwEjhpaDNnPp
EGTou29OfC8ZcIGFUukVLRejLsVlokanJG4gsV9rOrB8
`protect end_protected
