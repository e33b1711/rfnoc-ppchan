`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CO4puAAk5BNPAa/Oms25HA7E/H5O0lPj+5iJbl10S4OFe7/5viAjwlhzDI2aSH7TzijU+HjXjHio
bVoS1ymqKw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PNI5o2ObtSeUnDpWb6UmdcJVKwr9420KjKjTqEQeLfL/MNWFjLq2j3aV0odhIQJUw/JEaSnDEGWQ
oIfozlsXQyHrG0gKq+Zwl8Hx77BNYDxCSAY74t9bOXH4ySAjBkmP5kehX65C5OeSi9JEGzeRag5F
XIU1Dl6YiheDYTcwTe8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JS9KOAl0Ojsd20oZ5WD5EjGuNyzQrFjThms5dHYLgv1rBND2C4dQO2rdI8ToaWkQqnDBi7yw5DYE
ek41LuvyTGjhL729LTc6neZMfMpCzDKJkCiwTyAfVBJ22eP8JbrfxC63Egg1pdmctq5QvG5g+6JH
rpwYQHAo/B0lW1uY82siNqmFFU8nc9LK6vptKbH6XGtRsBAXaL9Shd1YUyUBHVXJ//U4xdIm3fkY
/qKR8alfD4mUjbKbE93dW7E4IJqSXWrpEkrL/ntUldqmdw8Xq9sHSYzVdteUGQCf8k4N0AmFibGC
RO2BJzt53XK5WXLRJ1zu9Pdqvb81j29jvdMQzQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jN/tdECHvKBiquY+uHEaeXmgr/LsBQSXlXkPeYbTzsaPKp3A+7a4j1fRKThKkI8e3mKdElL3llIu
/hlLmKLZYy4E+s0o1h7uLtDlFWU0yhwhnYl+4FN6Who4TLBZV8a/iylt8ASDKrhAGST6f42snM7x
LNzCA7H6sQ8KVGNds4E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bx+6IVe8tyEHkCXOCHEEl+1gu/INW4KDYqt87jjUgef7/prHiJLB0y/ASiMPcdrygLXZCainEmHQ
xiJW8SENDsmtle55onC2nitZvKqCYk0NL/TuUentDi4tONU8UDp8fWBHjxFXJVoIe6HpSxaZSWw2
A2bdJH6Kypw2C8fCohpuLwlrSilm9Lhokh/OCps1KU1yCsyALijhEJTqcHilHji5mbBHCuno9cbC
gX+6o23f9GSJeWwdni6odRu0tCIcx0/Q0P7mkOCQ1uTn6MmBJYxh4ucC7MvzVEUCsCSOXcffip9M
+aMa1LSSuyA+Iy4mhZX6d7hkf5lRgAb86CAxvA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JJGwqlu+ggMzoieNxa+v6vZaWBufNJ0QgHm+lgKECHPI3gzK7ORr5Y1R++Q1gE3F84vPIi7NxRlx
piVCdVHo6sO2PXolqvS14p3UTxW+rYskP4xPrLu3lonWRYrfunocAQff70SR7UbFfbkQCV+cOGQV
Jwa9pgPoTkYHyjhg02xm9k199V0mgIQl3GOCssx7ZjAlt3JjJwKR5BFVcNoyt/qEpWrKLM+BjnxU
YGZz/Yuikof8VGAFu/9zNQj4AgsKV5AK0XfcydwaaPGazCanWhuGc5ieoEIsT/O4+uDz8noYKOKJ
F7Q4zrJdOClWlbkFOLV51ULCq2PrFzKLje6W9g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13840)
`protect data_block
SkgO+InaDGOuL1LvRTi/yZe3MM4P36muNKNsJlNy6BGKEp88vjkm0oWR2iX2zeuU9p2YhJYBp3+E
cCkG0Ml65GVEebAfoKzhqXrB1Ss/KDtJqOQG0yiLJJKtjmlKXIlU5OYXQNggJxbUGBe390RM6Nsf
d3CIpWF6XNScoblUf60ZpI6ZbyYrJnwRxs/0DHrfFOcVULv36vcs1DXQ+tweLwSYFc5iwc6guUI6
UoaC0YC4JqX/tWber6Vif817XoxWlgb2ujg6AwriN3uvm6fCKfpxgDzyEVRLM+40qO+UVmDoBIRB
/Ws2fFq0sRZOzPu2ltnoI+vAPA8qt+VeNAwObm/aHHxn1nU/YmchaDGU2+wDcm1sCmHeK3oyhINQ
0vKDtGx6HzD40k7gpobACmv5R3UDoF7D8JD17zI8TCRdyN4EU2OYu3Mm3eD3ZzZBQBgCIjHWDdEe
UnVgYzDzB/AUXrLebW73EYPuMLt1Mer7xLxavgCu7GK6dEmwSU6DqPQaCc0u+k3nD2lK45urKBdh
kijgfSCDB/nyOIxlN2T6fIpbi6P8G6jMTqu7s6icnmVMPFBDEIFxObfPjHwPXzORtFnjz9ZZ7Zuc
M5cmGUmkZILFlH25NALUfYdqoOzKx+gmlnecvRwarP54485EI7aUgndFyGuRbk1SpggtdAIpmxrR
ZCCX7dm/stoULJZB8m2sVr9+B15i9NkKfyMueiRX1/DoUvcH3K2c5yrX8Ui6OyGBLbd1pqYZg4ah
hnx0xjgGNP+3SG3HQpkYRY7DT0cnL12Cye6vDJBJRTKYR4QclAZN1jeQn5oOCGYjhz8+be0ycjUm
qx8T6Ih+HKurOxeDAG2gUsV86GcOrX4kgIqHmipwv0WZScDgRvdteiv8CcdW+1CkEgBX5AppfGcG
2KgCdrxGaay7U3CsdRj60OrhFSBEJpTKsM9jU2Z0EYl1ORlX6lrIneJI2akyM6A+Ja3wiJAqxJiW
EzjgAFRVZQJUhqmQEwKWDyoB60RzF2jhjlWNlDv/R4aNgSu4jc5PTTst2Gxn7pKy5Jiv89U+xVom
9ALHgU4aPZOhJvfvI4RIG9sdE1xjwKsyx/MSEENy7GcO3vHgrhgJRP7ZEtKyX431b084SzCT38Ms
+IEZVA55cncHakzV3s0V62nDjVyCF4kRZPXUjG1p4X8PV3Psdp/6SF57SQsDeVqdLMhSnO9h6hjq
Jk6LcYqI0wGVTOcrpzR9L8ALsdgZdH5f4q3A9zDPIURT7xp/2T1xl4t45t6s42DswvCoPywdmIoJ
OlH445Q6zamAmeWBk6PwklKJ93rFtZ1xkw29TGRcTKo/6EwO7l8e4LnBmnBkvfCHSPl3KH/TwP1V
YuENNTjBJ7BKdYi+ouaPcQhxjfeIQZ3OyVXpZPkI4umxwUrsi5k0bl5A1wDfeJPh3wZNcwOPEOp2
G1lrN4ttOyM44YpJGXJhwfQL2Hxvs/lgdw0XHx7KFWG1erlnb5zNhsve5rcbE2XaYPjGTH0c6UaH
bteqSSlmcwd1ZyBUo0QTtIyXEUQcnL0MWZWbjemVmmSYVmoYHIp0mkN7aSTgwZg0zGlIb+KeGdRL
MNX3BKKQltqke8XRp6YDHNX+o5lrnlVWKLpOT6OWxh7U5IhfYklg2WNcTnECwXZNL62APqKg9ePH
P8S2BfIJEBTAT0s12ykwvLbGSigLti4B3VdINP3r2LZWfzlRk4ORSB2aqQm9ic+uLsmt14AdcpLO
SAKQBZCc0QgTG8Lv2L7bkT5y6qqjyeUCtB0r3yNt6UgDhbH9+MKvi8xnZOxVm+ENEUMW9XKBTMyf
zunGLZaQx51EBacT51jIIQl1t7AGXy0rvAD5v9rAEbW8W70nAW2n+/2s6/u9j8LCqN5FNodIQbmK
IRHb42ZxYM7X3uQwaVMrIr+fQNCKOtnY9hBOwkutIRzyKvB5dHCEVc8n6kGxN5LoAbgH/Yv6Z1zp
TMnPoTM08sz9aCr8EiguAH9Qn78lqZ3j8Yi6XdNIYw7LMpkoj1lLCqe4gkc7OaeH1UlAmpvWp+W7
fzLiYk7fv5z6YoYNKP2/QVksg+xZ3HddBnNkf8Dd1V9//PFwisvHkEcQEvg2RMw7nG1EZAB3AQ2Y
OUFzcjl9AfbXCKgHm130dvV8MsJIl8dizVlQxIEnsnKQ09jzgYblNOSWiVVnT5OzP8xE2EzXxcY+
wwHoqnC7blp2jeDO2SSDYXEDMMAqzJ8hxrFR9soaicri3LRf3T3cF/OzccrniTw8+ek5h8NVvqtz
oLz08OUdxepEyhQF7TV0g9NE8i3S3WuYrw9TNzVu9BQwM2rm0zSQELc1yIilJo3Ktkk6vpHTc808
Jt3l9ieTz4E3Nx97/aDbFShAEkAZ4U4l0l+rQQlQjywmM6GfuIOmw9KWAoETcYrkA/sPZgvpB1eL
8E2DZtkk/jPN+fSC+nQXiLMWfCrL+wEviVQB+5jKGeUYB/QehCXa7VgVPnJ89BEK+KLZbvqyuCtP
v/Xk6yRmMVGkDsIMdpLHAMR0OmBxu7CX2FUbQ2SinkDj0AC3fXK/yH17QOKiW8E3cZzDXGgzPi78
RjcsVnUeHTWFmWpe5/BaBRxG0IKhnjlMg2EyOFQdi4B1VbQB36IRhncZz+r5JyHw93ozoZtofZVA
Men/PRtJ0/D5qgYULqmkSuTbzlzQxVAniqs5iU1M3x3rg8EkCxsyOgTumflVBWZDRFqza/9/408k
f5UriVdZHTrZNrK0fbmzHGNFn0h7uuH3/tamVDXlJePnWLe0OXPnX5m0A2QFAcVQak004o93PMIg
XHb+q5SnHUwaAPH2e/T+mZNQ8M1JaKWhYLdHKifdvF0oEfnQMTt9ezVRWl/ZWqGbgS3KWRMCXHng
qD1oiEhOhpeswkR095UP7ZSFZJYzyTRXgcL4HW3TG8GFYrhvd0QLtCZ0ajFFGan96JS4IUcNyL/8
J03IKttIuAotwhQ72rePsXiSZQ40MB7J9GaSB64k1x6U7+MA5re4w2VzVlV9wTt46gpz6PKqGTaY
NRZfkhB48g8TA7oKDhzxGQQmfEKwK9i58GX/U2Bivju4JLInX36fEdIUFI7GysQyLaKzAqVDKDDp
5Uc6WtOSmZx49He0KR4ldStpM5i5VSkmyLIsh7csTj8NCJd9S3ZKHZSI9CXX79JhU00yaTr0H2b7
f3A+7Y0af5OMr9404zoOFn+Rglu4/4R020KY/77RP+EMIHumZpeXEHaaDkeYRL6c+iP/H30F06FY
YUTjQIVug+otXLJoXD2MRJY2+2wcAQElG8ghpsAFgdSQcF19YvhlIjUksup9CdqkRpdXzv2z99iy
MqWFPUhOFIXrrWbYjl3x3G2CDnPrjmTV5QWvw9dNBaRUvKVPusc5IzIcPk4456IVvZAVzxV6vdRA
tTFbK5Fx+UtfGOuSyNAZAzpWeHVfz9JvSj1jGazcsvOvTz8kVR5jf/jU8srd6eUUl0r+2B8SaCNV
Oj0ZGJwTqp36fw1TXZeHRrvgqohG3LBPGYbxjP9QNUIFyttbM2uFCd0poKBpg0WsSm6tIc77SIf+
9OeuLOmNCGnBTOCf9vEoRDEt3FVPZo+rNKubMeIhz3M5pbQSAS1OdaAGMR4+DhOLwUo3JysXrkub
u2CrtDXb4RLlvxSACg5ul1zBKxDSn+4RSGwHWLh8X3n/UePv8S/tH4vdbrjJho7mvoQU7qvcU1ST
cw9AfjL5JFdqXDV3ZFORHup1CbLhTgIVLynjaDmbzXqFMcZZYAy2qhnuldnXZA2r8o/Xww/znAXV
bibz9sx02GNNsY6DJ9Lji6KNlCKRyGp6kiQ4KA/UO3NF/CJofOCmOubDV7GiVxzRAvY15paLMbx2
Kiie9Rac6wPjnGw83SJbjEWld01GuS8VijCwTHyf0or2vUljJM4S5gxyDaLgFTwz4x8akiX0ic/P
AXP02s1fX8C55aGlmzfMdqH8pDJ9g15WbClPNH/Y0Csrzh+VO3g47RLBneSu4A06ejUvZCrh8U7C
/2taqPX3HqvPctk5oyCBZCSEAY+xSl+matvMrb4KyqOAsCLg83ZsE/XWDwgTfnQDp5ZxmUI5ce5n
w/QKdMzVpITVx0Jqce4iijflv62BSgeO6n31vUEfRTgmLoAi7uYaGgXIzHoQTKV5Z9bygQqaUkUz
fso/s802ie49O0ZfzOZTay5Devrbgea9yI1q5mI/E1igyEGKgMviKgkEaffNqE+s8jdjAQ/wvep5
nA9co4TQoEqbvbe3ck57vNR9hbSOTbquG9/+CBXEeO7jR5xkcOQLCSWVy5yJxGHzd9OS3uRIXxzH
OaQvGlxiUZsgCuMePGnSU2C3e3liSXER+E/T1u5WBhAgIXTFyYWgDvy5h+Sz+/KSLbn3cTP90jBV
JHDjBd1SBM81UTsLoeRbcwys5iByTWmRfdqtmiDI0Lwk4lA13LZ4tDI038BocAoPr6tStUf5UY4/
Z2edIGSInOYU5LDCg6LIW//OSSBJVYcLwr4WOAfXUUECVBV9KrJXQRTiDLHDBsWVKadTAtiAmV+y
ocIhVpXDI4G4GWnSmtPFN0V7jo6nNhjVGXECX21RQWYlAOwLGwKEZ/3tTq9m5y806Fr4QBuF+V9p
fIktYJ0NM6rH+HBvZhF/iUQ9BOJ6vlOpSr2x6fdEPyzy04O4n1yp/I0dDWyICoH7d/0PZElUriC1
SBIGRJaUm7m/YhJS/GFrOGOyCDE/6mP4ve57trKdqFKsV7ml8QxmOtCEF64YTkcoWLszVB7FzuZn
3HOSm6Obc/DPFaTROT88TufEZ+DTJ4jYkd0hzuCpNhrCCgxREuu2uh7uAdGe+77Sxqz/QzKzwjbU
p+Y5N1Vv1pQa3bkExqyrEUQyj/PujtNdb/HJ8+SrwiB3vcDCbk5kN6dwwXKrum9udAwZP1iQx/ar
1spGK5ktsiqdfA0v78LTp5EQeePtcV6arGe9Cw/SLZtpWZ8btCM68df2yCD7w0wC1mQa3Ryj5fHs
yJifOmcktxEGrz7E4peZLBLRFITaTSXJh15L1izTtodSDLDACHd3Tukls4AJlnYLLnYOKimvdial
vS/7Lw3WYAGa7nqMGfS4Puelr/C9TmyNgHRGYnq+UYGYkRg0iNSQrC4PCUJqT53ITp+05brnGXbH
6CRqBieeuQWb6ymUvKO2q8NWWOA+I97XWyeIPrvq4T/Llrd+36F1Q4YOspJ8J+r07TV4BxxOk+LB
qjo4LR/S9lcxxpc29P4ZcQZTuZ1LprdILmgI/qj2U/hBroSLS/PwD2KdQ+ZujR+NxqM8Jn/1jXSR
xYn9OZhOxdRpFhZAQeXECu6O68+2zCbONtomqD/6sLTo3MjQRX2zs9QHtVE3SV62hbEximnBpSgj
X0mgcBtf3XYH168r9GVIA6ZL126SWjAQByOzpL3UuG6V/QfCMpr3Jeiyfkz6IxcxINnQ0HA1nOX/
j/4n8BlHlcOmrhHNH3VOU2SHv6ASn1kQhma9KO051OKNv5nP434l54ypttbHi3gMeAXnhaGySlfr
lxI3lZaoCXueLcfFJTuSH1YGiDIa0eJ4x/mU4eZE/c/WQPM/v6lH+a6n+Tf9hUPVfM64SPAsKM2z
lODyR4we3kHZ/xum03uhZjZdbWTtjmGLv8I4p8qkQes1rMJSs5uoSYIlp+skuOL/3b4FTvAByL1l
CNRTPj3YVN/9o0EzMDl09EpGpWlmrHaaBADtKktzWiYPo7NLJqBrTL91ruli6TnXMeBP+/X8WaO4
1mPFJ+McNu+oEagoFpdu2CEZ5YRitwoGFNixA3QxtkB6yu0SiJbFRSB/VjwHWhA7SlghSR1L8A4Y
3H9+cKnQschHC9yOeLOfb14qLe9/kUhcA0iWAzAy119jYRnGTuixHiUcj6Duh8LKQaCMPyqd9M1n
afpR0wgwWAvqehsQGAe+jwIm9mboRYXgYxpmAFNhDgbm65mWNn0idvAwv+xVCgmTDJ9ODNiaG9I5
Xj4MGMAy6pgokQByanzG0PQ+uO/a/DjpkYcZeymwPyVEH/Reixw0XUqjPTdITmzhZ7GqUTgugW8k
V89falwNE+zuR4E+HH3OQz3N24vmgYBQjfitN7cpJgV8Go44PQImlLxywG2VaUqE4p2gP1bwGh9t
lmKs0sTRYtV0A7X8/WW4ukJ3WQnUvhY8zKG6HOgiFBLkSYNNXHV8fRTuY0FV/ly6J2qprKqkWYqF
9zrRueZs+l+CbhXgbLs4VFrkUubCw+fwCYKAISMu/w63mMSeyGRZ+rWze9a1y2VLX/eKOvJDsSWJ
xlfzfB7x8ebbTsV/6jsUOQmnArCFsWhyuDHmnEmV1DFQ4bZjIFRXEyZLs00Og+UzVw3CCPyGbb4A
U/d8S7H5Ybg6rsywXiLzuEBrc4ZW7CemSFNWNCnXDNxHQ6XHBpww/5o2rwkyq5j6rsB19o2Wp2xA
BWs6rV1nl59J6OKXew++IMLLtc+5KC3OOP653ZPeurK0oE7Fe+fsgkJcWgOU/0LW1J25V08mPqMX
1Y6z/C5qCztMard+Tk57QX1EuDC9z/MH/NG1R77d0vPf+LmcXNvVP5jM8R1i2LydEPhDbReurE3H
BZiygvntDZcAt+dvKdmeGAOg3IpYBn84EuPxcGNzDwna5vme0JhIe3RJc0/3nCBnXrNELN5nW+k6
6Bw9KwcBobs4JV6vDC2kQ4HzY0zA8fgY4qJE44IlmranQ6sD6L2PW1a0C23pWPMHozO8RvjygFkm
brBm4ssfsgBH0D/1zireZgDXyRX4vtKeARVVNvAdS6sZwOF544FLmpxnvqyc/B56mQKObYT4qJ2S
WO0mtcQSqswdwpftIEH0MXRlmpN1YxoljCifUfMt8TibAZ8WbpIzzjZ7Fg5XMJBCQocEkHeA/bWY
nGvGY1dz3dkORBSd9PoXyS3cmKBTlvvoyiC/i9wZM9JISAOiTpyTgdFVMQVtNtgXJpve/FjCIboB
RSCpOlnZfkDCQg/AbObt9YINCZYKi6fuaCEZr3xwBV71yhvbxmRvNT0G/7jTzKCwVMEuW9Djh0bH
N5fEbHbL8jL/fdtH+3vpq3xgcto39A9GDpCMncGbpAfmilz7GmzmlSJ9ay4Qy0LEfUuFSmN/jFLF
my/svI47UiY6wHHgrCXHwCY5Bu/8tVIBhsYi2+tNQuCQawIPoLnHzZhrgxxBQIDXd0WcfCPaovHW
dqgz6zEJAsJq2YBlHyvo5g9c7hEMO4CbRWAJTJ8UWrddKWbdOVpnWXg/AhbeK/OBkJxfn14jYn+e
4qCvkBtK2OPMNqTJNDtpsPa9LjNzfvWGA2IQDAb2AyRrd2kaQQHO1w4xpguJqOK+ZZZ47HSnR2KM
QZ8V0NppGWphEhBC2d7j/lp0Tppnr9m2zEvrM4A7VZr/yOqgI2p5ZmdBGDl2CmZIFpcEJa+Iml67
FpP0huVd2Me3+ZGyQuNlevv9ocr08t9Atlu09ZP1mC+N9paBKRuWll59c5a9S11M7d33FGbA5H4F
6rZU96PuH7pK14WBTjhmcDvJ2Lqp58a4AbM25eeBp+3IX9/E5p6mx/WaH4brq6xVQdN2bC1B0HQx
KX0dXN+Fja6NE2lbqNPvWMC0B6dLxwKOS4zVVOVCVOsNOsNqldWahcTsMfMF56OGL1N45aQGlMjK
cuTX1WmmAptTGMrIvRhP2HjofWRuYRTJehTIvJezxMG/ESGI3r71MNweVL7jtF0OW5ThRGaqRNBC
u7/lctMd4PN8G/d1Z8I3hyKzk8UicrJMRMBkZJ9eBe/xRt+jCQXf2Lk6iOKGYrzvLN+/1Hd3Ds50
QnaAgfEfR63hfW+jWb2suxnMM5CJ6GWssXRbMfyBNXMxIa33NeAWnXPbsmvgK2bnpOis3GIuSdRn
7OMNZx9qaYngvsx4RghB1pVQGdEVzqGpyJBPt7P8isxNRoBpT72aVj1B3v2CRVkbgdcQBJi6kU4y
OaekUeAofSGEHZNimfytDOoa/ch9WpyUpYQttrwXxqg+qKwqW0jg9PqdmxZm3eND0FnUPO7t5J6l
bs3FEfXQaR/SoJ6Fvml2bOH9FhjgJeKay+3i+LB5bNws7TAzVab7D/uh9Bl5Zes6gLvTiyw7U/PU
dFOQ3MVug7KRfdEcO7JI4gLdc5ktsesvnZ5W/kX6el9QtsCoUsEyDPq6ZJQZb5Cbp4lt+KiNP1LO
AZBUGVyudJx1+6nDEANyP5Ha5p0F0ekLHYiSwxaiqp7n1qMja06+rUgbdn27gJrXc9dr/N/sA7zS
VpWnljoDdaUO2GXkLrjajfWahhCBNdQUjTWDI/qCmMoDpAbuZS4BUi/n+m0cimTwjs9VgdF97eGq
tue+l0803LY+d1J1Mv+cEd3GaP/V4f0aFNo6dXf+232bLAYbMlI7mwHoZluvNFksBd2zZzZ4Y4fk
zJbs+2m3bfShxFSpckDfYtjVz8wg4sx7Asmop04OCTURmn35ZQ1iQixOnxRe4eymsvTjc28g7H32
4LamLtkLS5A1rsFcyyWFNRDvXZuKJJ4OcXwyHHjWSsWxCbb6Q/oBdPFrYlfWTyGrcWVL6CtVJXOp
70Mgsq6DPEYr19PJpTxslXu4xaHmL9ApBvN44QExzamkGGbk9VNM5IGQovJ9ob6uakbl407JXZZo
yLbGJGzt6HAKVw6JdMO7LboXRr/IQV5jgYQmSjpSxDJaGGhf0YbXComGI0bEfswVLBGjo28SlgDe
au9UZ4je5457/AOoJGsQDatsrBzA3bq9WxvGT0H6tGe1W/SF2fxuoLDUJ5KrXWCaHXnJJc6rnnwP
nZ5sRB4qGmMDVZ1fLEGWelH18PFgHaBKM2+OYkPMG35TBJ0It1Xz8ezRb0SYGa2C3hCqbnOIRx8Z
ACZEZnkQ1gXRckkqnIDSPzzlWn0f4WUHkkIwu84fkK0guEcBmZmNOIXId3q8NT7r3L4FDVTJhAdU
S1WdGMJxCovsnh0ZNSjPaIk4cnOuxbguHoL5/evK0/iv1inQTAlYGAHZHODEbQ8bDJ5DXeHB9/kk
qeNMyJjX2BAg3b4bRwpAVBns7/a9Gtylgc8zV8zCH+U3hTfmTriuMkHOU5IApwsES+WjZva/aOYw
xMhiK+G3OYDIvJS6yuTPB+jT+sb/Yenq0FtJEJzoq+UzQpAPpJQ4Jx/BcJkWgarlhPTV63+0+oez
64z7nZyUc7ooyvBSMZrEqR3g5q3Eedy2JvvRpBO3ktp5qOPhoL18y7yOHi17UPbNzKsbcvs/xVG9
WGuQvt9oj7ljVqVm0/GITnQhmWmzsETknRDxHwZtUTNLSnump7LPcriyxgl6PUNSv1VqxoQvOGLH
tXWTmYXcBa3mUZshCYkGNSgjnGP1vy5Ifb9Xt8Kn4Y3oAkjpA+PjN2vnaXE4VrPEajbccVOeW1+g
XSGaqRYNz1zpr0yMYBnQthIxxLJ/ZELPKXV7Tvou6nEFvxYoQ7nzELVjv5ZihHvypNk23g93AxsS
YFPWbdJaWBUEk83LSrnmcCmqp3e5wmvXzia6jAhpw1T0yONGHIBNZ5bf20JwRZnR/7qHwl65Xkwh
w2uPxwUvLlPACLShRrf6Q00CUPnRFqbBzL0AYfwhxGYFUBsE95cN/Rl9TQDD577cpAoxcp/tGbjY
a8+ZXjsqJzG18KfOIk0dMatvUzghINwGIA3uP4Bqmo/ZnRW98fBoKpq2qHvIcGWMzaubQezFl22F
SGpkctUTH3hzwC59XZLaI4XFfTB/1Sg/0Y2EroiK7ev6slPXgqItD+AGlQdmGRiyp8Bd3gBulnOL
jwmECQqNqAeKexwdq+iDjrFfFVATbIwYCkmSOcDpVa9KyeJJfP4xQGYy08OfbnP1m885Y+zWorNP
SMcxf/p5l+C8SAiUt1yvC2fesIXs4gJZHRoSNZHbFJKv8e61MrOflfxnuTe9Lz2dZUc2ypTcXROx
5cA0UJwGhfpfuHXt5Jm1IT/veFDc9zDrOg4xqcWEPDizggTn74NmNIaMoRrXIDBjLBSK16Lxmtbl
tHeVQmBQpCdEUvUqysfyszBO8y+80nzk/80J9UTpjb1gGXzTsH3pu/Y/jyzO0cv/HdVqH6utwYzb
oP3PWRJNC3Rs+oNYIqNQeK/tINRu8xDJYxeFuGEbk4HaGV5AlgblTyRmMrsriK9Q+9JxZw3tZO2F
SkF1UUZA926ZEZxE96/E2tuZ93I79j5cYs+uSjEAPUiEeqfNqSfi0aaGlH99vwAjtg18n5E3jkrn
IMgzUhWntMheY67Zaj/+/uT0RRVwRxL7c4fpwIhQLv1dkwPcqDGUiUjtS9pod8hR2CoKBQHNkVSu
RCB9LxqgIW4FmNOLJRxGJb15u5pLEmafI8D/V0apYYRP1RgXvQKDfejVwvDUCAiTVlN+9U55cc3T
Kp7ZqW3jEiJk6WTuOem357THH0rT972dSjjqa72UwUeLk6Ei1hv5HEtiQdIbrI2AGTzrMKsrQfVz
eCyBbgK2mhitIwlCV7wm9KMUWvWEMmSNQqXUTv6d3lTcqRvD15/58cDIzVuBbKNx1s+Cl9UtRmv9
vApZAqG82klfsiQLGUMnUCPhDRer7EjHzSUomoQKJClCtSFwW2hblAD5Ra2XKgYKpQaW6kalWaOn
jblQWldNDyCcZuubodCOMaG4O66gZClV5CHJZcDxMUMGiP/vF43N2m8GdWEMhZxRjDHHYZxwPexO
6wQTV1SqD2FhAQIGYsGyxMKszniNMKEegbzjDNidHEK/1pMfsVPfOeK9hQvxPdonh2D1rihDR7Ps
r3nAviuZBtns8OBSJjT/JRymspkNTwaJgBYJrSch16+KylUZmRX6Zmzca9LcXmarx3Ur7iTnUvi1
8MlmHSRClEBUNCJFo7aHYc4S6W6YlOcLkEiq7PPuzRbe+iuMj3/bYiEIF8pHQHAORh6t9PneISTZ
Xz5lhDhjRVL7aQSwmrsFgCJyDsPsB50dwDpefrqGxw2KqGA7ypIX9hLYH0l+yXFozmQC+WG6lGtB
xFyir2KP/4/+NwiWA+9YzZClWmuhyyZwMnVkqraAKn4MsPzeUnpBzaVRPNx0GoqkvZxdVg1QvBzf
HOflwS0H/jSeWWMMk1PR7Np+J2E1kcLn5QPv6Ge3As4nLr8LgNcwnnLVXcCgvQDaaxfg5llP2/vU
Deh90FhQD5dinwE0xB+Mt3SIGHJN+bCHildL8mu0/xeAQDV+OG4T43/8hdvAId3Pa0quXWRQru/e
H4lpGy2ukJvJsF2wME/vhEHx2/crD/Vo6UzJihEM3Z8iGka4o6XRSCH4m0sniY/EoICcdZTl21VX
Afdgu4cKCKb51LdVrGxSWBNMgLRmLIxJviSUkCyX5gL9zDUQ485XvubNkF4AkQC7jSjOXqsU/WoZ
+fcYnZ/ucX0IrCNmK2A+HbQ/kfeP1vbr7SBlGtoG4hR4o1twAQ0Zbp/45qIQK3dg8lvv+t2arneK
Bgt/sAN30JzpwqgxltwVWR1cQPwsQMjG7hekCYb6D5dQ/OKykaTi9EgxfK3ODdlNGeVJc5ZbWe6w
BSLxn1SEcqL9i6nO8wchXFgzPaLZS5ldvYzM83PI6VKbCk6zZwf9cbbDKF5AHZJ7NHsyrwBhAXGV
71+O17ZE5EedJ0FD1cTHexLcpesmV/vKAI9UO1z7Itdg6xaptLpPo+HqXVEZAIAPtrglg16IeWMK
1zRB4mI272FapbCD/wgupxaKh+3xjganQ9S/bi4ajRVm9nO6ULUDe/1Zf/D6VeuAkuWI7eBtNT93
ZuWpdOtObklBWiXkyREOuITdgve7OdIscNXfjFxblWvpmQ1JdNH/g2+Ncda8ngGSpEct/ESB/fRs
SOn4YiX5G9cPlsucZRzfXslSdNtFtPkpMPj2FXw23DIHUx59bSMZC2ecUU8QmZ0PjyxB8dxrkJor
R86R+5E8vmKi8HQzHMyqaqjvvvBxEIwblVIuPim5IRAL/60YkQE4GjTgpiGI3Qf01oqlXjFM3gVJ
1f+rkYE7hPhD31Zh68eyZudXCPtGk132+58ABHqCBJEl6PSFuoh+w3YY3wvUKVW95SJf3Q32RZfo
hBaf7lYECIsipulxrespr2jU92bcATLnTbDQrR5BmjRLMWjcPcfZdSd2NNeBp+5n7HwL4LyXxg/p
2rgQCA6rc3ixIVyT12CYp+ljJ+nNsuTYU7VKyxvoxTQcgAYdB4jw2Q5Tq1f72rZHECMOFF506uTj
eEWy+ZXTsTsTQPdvGR+0RH75buhcmCknO2EJe/p5qoD9AQ+9pw/X3ThtCBzCjRcO7eFoR8v9bUtZ
Mk1QJjLzV1ncUhHGNHql6gwoguxd6FuHvIdn9JJa1eVyRgmyg5tFJMXNDcjWuFUyjSzasO4PpL/0
JCjL2XKUpxbMu+I0o7ALvyptJpHBX7APy4Vnta2qiMTxdtXk3qMkBGXccW94FoYAvaC+4qiYk4is
R+4qno2zFYi/7YnGaw+8bdXcU1BodIfr60qYqg14x23qQQGunaHjGBuRiVsr2auB+Y92iSQvWKR6
930uecvnQkc9sk/EkMCjFV3bQmBLTvESPUzCyRkm3cMoBMgKgdeiZQLyM+eCn+/XKZ75mGbzAoHb
NCFohJN3j+5tUqNdLaheXVuscStrO+K7ba46FQkY9bNZp7QiGK28xVgv7ruxAop2VDz8zbcTn3eW
fPxRC0x9fpT5CW7+3m4AeF9JhMXpDr6amyOzumBeNLDkkD7GR6AtuVjOGA3yegSFlDPlXYgaNFKM
B7qYOTdINRyYMhPLDEYtclydrD92tdqyS4SXDFntZ0QH3wBYNEqyt07CVaDTYJax7sFoA+uMn23M
9ACMNBrui9g3/Bxc07eeAC9NaR9ilVTV62kSFZzqGcIRy9W1UlgJrNXXEUnRiaen9lXYpUtRHlVL
Kk6NNAGoQM/b1nKvGpvm86Du0/yLP0T+fI05/e8DmXvXhdR0VgrbckyvOHoxCZKNX6dTkivGJO1H
OikFgs4o8pwrZsp8vO0YIaOyIXVP2YTBUf/PrPp3zluGSjWgnywzQRbK+K9tKxwJy3S45mQfbWZA
8q10HaNSX3vljkfYyymc5d5EGdb6ddAmzD1GzfzCXsPM3kN4RNjVf9xsnAnHHPxPth4jmuPGBLX5
Q7ZLkIDombvMmarK8QasCnXAR++YAriaGlKd6u9qQv1hyxs8EuIbd2b4MdpbG6x+gEbmclLznFYT
29Rky2lQL3NepWuKNq1rYgDXRhHIFq65VrdmxmwgXgvCDKzN1I+WULJvheMoO1F2FcpTrCkcsjDI
SZxyx2fqt7MUDBX/J0PFvaYqEkR9YnLRFZG3Snct8wkU1jivmJEBxrr8OKjOlUI2UnG9cd8PtgeY
aDPJI92uZeu0rP2ZfzPYa3y6cdCRMcO489jJu8qzLrY9i6bGiIMFPl0GeWqv1FNKmsEUjIOxvaQk
GbXtYV1Zi19EXx8FBCv0u0GbK0kyFzNZ6vX6S2uOerLrGF9b7qDjDaPXwbkd8XeSJAMi89q4dBq2
eaE2dzyfwRWCyM34go+B39WdStQCdLgddaFAXkPOn1cFwZidtQYzWnvtf8Qz2RM2ojMmxqv9Yq9b
3nGk+MosEMqoLAZbvuAi+r2amJbfF3G0PvYKB5g6eHG0y0NxjUPzuYhU8dSV1EHPERctA8dI2iyd
+D6LHPZnL3o4b9vF2aMIicK+zx34PnRIhwGCS00ec2lnxvrSBnJmZD8TTBafFZjE5ZLY9V9YGAl9
fVvYU0Xj6MFpMoYTJdr2k9vZgZBrrC76fdFn7eC6jex8FeNFrl0Z2TvCzOi/+c3GkrmmsAaJlqUO
XutXpvVIOoTUurIL31XQvQs2aIyqYjTAJD6MSzL3GHUTrnA184n/vv8dfMAbtGQzQFcoFvKdVQvb
noMBPBaBC5lIz0mFhm/sXPHNo1SH4i2BWZfF5NmjztL0ZS+ie3R76CO8QCQ1zeyRl8zZ+8yfhKhg
rnIWLgssCMOx23HY23bNz1R8zY4zuIshvWEReKflSONczlYbh6QsaHXa9GGIbHzu1/yqv+C3+u7C
AxvHY454mp4q5wYmzFCo+9oI68eX3XtggGqfctbLqc6aIT9YTz8hpGpQVcMWj0jERYmyEYoKRR/J
CIUyrtcNy6isBxOnK9eandEifWfVSnmCFa1UQLmTz8nSVyfcdkAIKq4iz+Y3IzlTuoEqZUCV3XrC
5Kidsk9ZlduvNxPIyvccBCYx8BThHD4UaRggs+rVhVoEDowy/7HcC6xnmFud79iic2bcbxJhuGN0
6F29hXWldMCGmeTyLIx4ciWR7aXQst34D4FSB1CxRJaq07sy3LtdiYMjtmUP27hIjq5DgMlkIwo+
qzUhsWif6vzhLCP0p4bV+QBQeg24Du3pMJmJvInY9yWw6/6gy/toIylHkf60h1pDAe5Roi7VozjH
6BPucClvaJUS84SnPFnbxd9v0KOjakWZJTH2vo81FwhHfcP2Ar7jT8QRg1/7iw5NmPHq01CBAwSn
CClggVTi4h7oqezhIpK6otsltboY3QVbBuE2/JdE3XkoGnvTItFQe/AQWlh6IUHweBXBDPQvQO+M
ToSmP4M3Q0XAOXp0d1DwaK35ym3hj6ZnfbkYfB6WgQrkR0l6wWe+lW/tGjS4oXjVjlp8syESmM2/
oMAn1s0ShqXF+xdRSc8LqReMsAVBm0pLag9ykf5iGI1rg7cPms5cJKEKm8wkf1/A3m1b3I7DOoGP
lLe7gW63iswbQnOjnLH5hi2jrJSuecjOYYgV81MD7WPypnpAupi7y+oqkQ9GT6lSAswPOCEWz8vp
6FdXA0D/uX5PngdLAdAniRN8OeD8UfxibG6vM0RzezLRwkjJGcYriQnUqADS2gAOMGM2OIirBBuL
BrLcFxjqyL+v0yfWNkSal0tL7pDRrK/TGnV6pXnUW6pZDPSt5jBqDkszIjGFSRrVvEZg1scWqhQJ
02+4f6mH2Y36wn7gj89MvyIXmMqikhHOuShbx98a3lLiAR/Yub9o/j4tn97yIyKq7QXsglbcIe2k
PYzZQRMxhjYBwBdXwYy8cbOa3k77GLcHtv9X/mpJqRbaHD86YAKQWqH/k2UsT5EwWXacgZNbZ1mo
rr8RH6DvgoKpY2UZr7zqdJI7pE0qMkgn0/3z7cuEjZ8ZZwZRRU+vuqgrtToAXzeNsay5PUU0jV29
syQeTBSBXoWtJPQz3RrAPSC1lu5Emw7F9dc2b64YoIXbxNCGkA6yB6KGuDoAywVHzq6MvCZ8AxHW
fmNQpdhK6oPmB7LYisBm+etvnM241uH6QJLEeaExK5ezQrW7EHCm9N5MTEzVwWk1XjRq7cHUqIAj
8CnbEEOnuBYooA1Bp1wdakuD/j0aRL7lov2RUwRZGF3m5kP7SmZZHiEQgmXNxV6R4bROYkBkpWtO
iWg1i7fZmk2GF7n/fHbDfQ1lNKXxSYyLQ1MZw9XJ0QcuG3iqKX8vFWhBp2BI1Is9f2bAqGtg3o+q
KDPNhV2+Y+4IbALpqiUH4tAn7VSc8vXFzaGOGpKjLMmeiFfNyTiVouFYqSmjDGtz5KZ2Tj8ZleXu
OjLi4+fOjGtEWF3CcmfOMMGIG/AquM9ZKjvqZkH9yNvmQj3LYff3qmhXgzw7dLeWu0McHU3XnOIT
oXuuaFpjJoGHsgKoHEhshk56h1ugLplt/mt0qWK1bB3+CCfUlWz/QpGO6ULJzB5gSD99DAXf0WSn
hiNLuMS0FaCaZtoMREUJxGJzrb2h1lLfS6jceaVUyYfgzFjVjN4ygWzwehHhOBG8HTWX4DhhepXN
ocQKkvKJUt09mYZi8fbbV6NgkMTD40adSUcMDEAF67t3hmB+dyVgPPmvOgl5x5hVaRBnQFca1whY
VrrAJyo4mVAJI9JOmMHmjfKpOzQYm0MfdJrmZB/sehvz2TS+VrEnBoevplf8d4+UeD0HL+H0K0ms
XNwTqXWCxjOM+1faCtClZuiDIiQsjF3m7bfQjhfweFJvMHj3h4dq4sd8+N4p5i9UomQs4leQZoLV
Ao8UmxLGI5+LALdkwQSIFnut26xu3KjNvFEzZU+xEkCUsBWaD8vRVU17ImnA+FA33fzEK0Q6t23E
jYMSF+Ei7OvGPQYcs56I+KK2dPg2k+nw24IvwYrRE6m5Pi0Q4ulhdkJL+SYohIUp957ZxYxWPzg/
PReATfa//ObivhJnkNOdOALsFZgRkJjDsdJK06+NOVTyTV78V57Jc2hmblbjZ1ml3iGN0lMvh9N+
CszPUoktwtuDuI3JeGaiz6qAl8aYHu8qCpkKpjNQ8uU2scVWEo4hx4NLw49YASU6Kmih/rcgXNzq
s5TVW3NaiyBWoswnRl8FA4DtgHVGQYCJanSFwYGhGla6AtfOHiUpHQpjnNewpGMvM/QK8gkihQl6
exSNFViEeXxe+STa/6nh4ZoxkmdblJqSN9OyLG7vEDdqYLtJjGzn0e6Gsu3X3HgdlWTYEBhD/mq3
X6I1xM2Mn3EwHMzNCcnrUZn9iSTBRDG2nsnT64lXbZD4IH9fsSajZZT3GYrm74f23hmo6LVLXqxV
ngPkKlBowZpbL6EVm1QinBOCeM+NN8o5Zg/8ie7OamHgr/GszbFabz7qoHLm2HwYh2s1I84oV8J1
pt+CRs2AxMXxr4Kh13Gn7kZAUlhqU6NY4jV8S1gPW+T1cHRsp1j6IriIMBOpN+NRqNoWaiTpBZ+V
dg9oRezroH0m8IXQDh0YHByJg4JMsVlkGzNz5GGb6WJ1MUFKXfVX9LP82+WD+CnMHGBxKTKmrG4m
pQPUfZnYxprdi93zqgmz990O1cJxDPlPtJU6VmXY/OMvLy8zrWt0Z/MA/O7N6/foaWO41iULyq/c
EO3KTo3PyrsYKGKAUm1RGnifCrG45RxY5i4ACkXfA66pAVJ/i6eY7lGGrD/fiXECgYO6+1f/TAjX
9Gctpo8VQgyo1ex8rA/Tka+j5DEoavLlVp8o3dv1wBFlCw+7ohSXqBdJBqQQKe6+FxMd6KX73eUO
ab8LNtzDfUAp5Ie8tlbd91ZsIlefKrI4TOuW6zGRaTPPlBhEdbI9dpJeQxosAiZF26fPULh1rVON
mbsZDXd1JUts504fNbHyGj2zWzm1DJ+0SYJV2fV1tBBoh0NzP6FeT47yr/1PCI0nj7iqbxjIwHhS
8vXeTAvx0vS4r9Vtbqz3jSy5vh1Sgey/SiwYc5Fks2u9OX8MVteDpzKgmoab7c+XwtbdhR28eczi
DTj/jz0+BZ6dvYdtDUjXvPVXD83AFJoUZeW6SPtr4NFAsPDPq6RnOZtC8qX5ZSwR3w5pfHK0zJI2
J7K3Z/N7+1wruzRVvubZmle+LzKI+UQEldQ8xrBUhT78tPfMfoDZKNsZTjJCVzCfwzaQ3BGtfRSG
GkTYw+GhvmBjm98/KgWsrtTeysp5z0GqRH1Oy4CeKfxaS/DtAvSS5edeNrHh3Jnz0jeaBFy9nfgJ
kNS4LITVjKRnN4BdOhRkrt9UB/zmjmLQW1fptoTM4f7Pe9Q1BAmB2R3e9BDq8caSWCqS6glG3rtu
TcVTOjI38BE5mAvpD2xBZFRsbAm5PVKFuj1D4lO72CAhsgKXWFQ6d8VfJXkzCzcJ1XXrSFWxYIhc
rUDuwsNpT/ghI3dIhcB8CKpVzplSD+G3VMEumCHrpbzEM2V7XqRkPug6rxTguqO4GJw41mnJ1slk
XjJi8qtIptQ49yzmGfsYG7PFlUw+Z0urRNrqdvVoRJR0tB6ZrQAxAP7hr2PLPdtDJn7a5dcNqMtU
JRNsCNfuQMlFnAHtzzu9h6Klc1vNbMaAWiph3jJ2lvVXm5UmnnlvlUIEZabrONT0UmfYmp8UVOqi
VLEZQyAtoIwz8A+zhaES2EwhLWUcOvCDUTw9twGEGA0B4fUY9vGmgsSXPUF+I8kq63BgfGkRorcV
iEHY/rjko9yx4EMuujY1tRWpdhMxTlkrmTMkBaLQlXIVFRRCgtvO+PVg2TDAJtUEzE4GEaIVkcas
8jc57wcr/zkm665XvGFvGGDFaGL53FRM0382PloijTdEYVLbHBJ+6zOXoE8+uZ/sOpmI4TnF6vPV
MTkOtckYB1R7VqOKqExyf/Y5AALMtZLgy5CcgJJVbr8HOcalmjHvpCC2hMf4FU237+De5Vq16Hy/
iTmFNxENhsmKhX1xQRYBvZGRUvCWjFAUlhpsGJN0qofBnv9/G/SomTToB6S4RooWJ8zj5RrqkIiK
5OSblCutf+iIccyDQCE3hQFj+y8cz+Z9GjU2/erqDjGvtZA2XdSfWb6ZH4k2EH1HptUYc/bXYtw0
Rk2xMqRANlf4exBGDgpXdO2MsWCI0NgQUcF01zVmglPpyYuJQNTf4tqhqkJfbei6bnNN5xE5EkuH
5409VzHfRoFgU6m1vp7XNA7t5A39htmQr9VZrm0fB5nY7YYxKOAatzbP+crMmw==
`protect end_protected
