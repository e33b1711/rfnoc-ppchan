`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B9EdoYjgQSD9gDMqVua2zJVflRHus/LVjvgqriMNBVhHK/84/U2ioEKVQOwfFeXzEQ+lX+hFCLqk
IZ7jFFR3eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RhpaDjajcReMSslu2NKOwc2kbW/sae+dRFDHfVBTDCkPzbh3mSiP7TZOBqhKDGqTB6232MKVx7qP
ZBtzaagM5AWVdbRcklCBM/Kdvk2QRYet2hF/9C2MMh5T893aaMICNr83Nm8Vp+EZuwMrlQi9gn4g
ywBMUWKYky2UWYxF3K4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EMspBr3PE9iUGaTBx7AjQJAXSHmvP3RUIoqkvAbDE+yVNcZvKmwd5igMnbjWzn6mF2c0q5bTEPiV
SW2sgdg6e+BWLSQSGz4p9DMI+GfIfZaVwwQEDESBje7X4DTUoGoCTuJszgnSgaxHrTunK6Mskti9
6KrQ+39Cj86aIm/Se8nuNq0dyvAGREfF8mO1NUC0gTq7uy5v/YguCmfE/DQabE0hSg1HMsyBV/Es
GiQUjqTbeVVWXfqfBUzosAXVQKO0zqx58iAqNL7CvcGEpsb03lni7FDq7sA6yXUkDI0QOTEsrc65
s6ZtU7tJTAb29hQhoHqIjiGrJFezQoQSsaoiug==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b93sxpNwCcwf4KNpCEGGFkec9bpq/IxvjyBQsUyVkA9gs5+mZCPe1ZsIgPAcV3LuAs/hO5uF5ZZg
8XlLtMGUzLOqudI5PSmMsrYFDtN3zZH6HVVdrqx1SI+iWh7n9QVxAWi0Gb+MTGVlekns5jXfAoVc
3u3FT2heMRrTJpych9M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bXZyR3Gjk3qu1g2YuorAQnE8wshy1nalVGdBpmgUZ44y9It3o4HVFeQyueq4jESAF2Ey1VYIbvPD
74ozsPhX0ixRYVusT9MV8PD3YG6LdUBXI17bxA0LAUmItJloxWSXa+t223FfWE7eNn3+E2em1yes
DofEMqIUoCSM1VrQfdWQHWipV5VENa16uK/O6WvUpm9HCeZutIr06Cd4/jMLDVN4zK+BRg6PzYin
7YtmQvIO/IfyaTOOFuJMXbkqdaYK3LMmByLBTTcc+Ph+MSoPOSUz0iJ+rEyUD+vUc++9MXYxYO1R
d+2oGZu//gKeC/sSjsNzj/WkgVmTtfVW9cP/BA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AskrFrWXFM7AzCqlwzwplr3AKnGiwwGzSK4bMSSxCba2xMWeQ3z633VSAcApQXs38MGCxBDDSYbX
nUzKzPFlZpAxD4jtBhFZhYrE2rfiXck3GhW3dp69xEgpUQlfw8i4t1/+iPNzpGa99NBOV/7wTUca
GQByFwIqxvt3bKLQVKoSCzYzVgdmM4ESHX39oRKLp1CBheiJrFmXRi0x2ea1efHoG3nUywaxhQeI
YzkcGouUEqPqhgI3U2ijlo/YVImbNvFBcG++cJWa4jTlqPyGPe3ENw0VgoihgHcOmdTWUcL0cLlB
R50AncMkumkCzB0MXaTqW4ee/PyvqhHRlRf5Bg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94528)
`protect data_block
FfpFEXU99vgoUXkUYb+7PKBszorS0/TR/seXQrvGwzza08ztCz3ZkvJTJcWr1IzH5xQcmZhZI+iw
vz8NaSTKhWtBWYtChBgIO1MM2hJt+PsR5MX8XCwDVSjC2BwXH/RCRdkB0dJ+jraVuxCPnvc72ERr
L6N4+qx6XcRCrLAVvFbK3ArandQy9VxuzpLz3R8hzNn4ramIJ3iV0CNoriS8lgDvaSAMwbG64kHA
G9JikGO85mU8jNHlfkLRzYdg11uQLNZl8zi3f+6gflPTC3sbkl3Dwny9HzOI2NdL3qBILWfXUU5A
G84taEAb8LbPGHqv64XwgbC2yNs7aImHZaZdN7BdaWjN0fsHE/u7Pa3p0/JP0lvz/hPi7JpM/S5A
5DoSZhhW1YJZmGGTaZVdllXmE05SNnS1t8X/oFGlwKjBC50Ayj2DsMzAotGu4Apzuhz85EO83h5E
EcXEIXiU7RakBKC2+ixPc/lWpxom5XUf/M7NQvW5siPHGf8i2k0bV2xEBe9nJzYbbHW24+tGcj1S
sakr0FXxO8Gl0d37SGidF09SHDikQaGMUxAkaG5h3wx/5EzBzH7zn8aGon58Cl32Mn1aLYRTLMGu
jc+yZqQW26LdVB1zUB2Y0jLfGn7fORTaHE4exR04t5aBr1arnkC/Cl0LdqgECKhSuuDkcJv7J3J7
ublxLd5PVlNlJ84JKmAglOu829uGS3k4DqfTwKzsH9/xD8oJDust5dRoxE32IvroHlAf9HBNd6pt
+drZa7X6QzVxr3/iq5XP5HPTMKATWC8nqWdLqeGuUeCkkGqeEEojt28zXjMyTaf4CNmTT56BBuPf
s5FfrESFLHjoIZboefLcK4pdfOkDLuYntC4ysVFOfbScNtIvyv6DuSK9fqwlWl3P8reEu4pflvxo
hrgsq9r1bUFA6pK+09ASdjvA9cCoqQQm1NERK3R7ahKlD04U+lH0uqufidsa53kcNWY6/rzI9oIU
lxdS/xbF+EazsVgqx+XohSBUcCanY2vgOyHEBuRXwi73AN7WeZqWuZ0k1QuYDwSia+kfuLczlVQt
LXeRnTtac/6NYUa05/2etz2+mjDoCjZn9ThY4bqzzy/3kb2pOQY9oT3te9TVAI0zzluogoJjtPr9
d0f47boGSd8DiqdtWMIoJhyjk0e4WK1BaTL2FJfpRFd87fMdjKy2q7mt7bRb3x1tkyfL+8jutMe3
qR0o1KhVlyvGzEGp4G1VopuJdndlcfjXMhR964n1MTQS3CtDlraoTmrozW0+7Qc/BRQCmRbkTEFY
7vawIdsADaJk124yV4CbNbfO+x7Pw1s8mCIzPODAXgVh+CJKw7Lh5GSc2JG4J0Ge8UQ/UTChwhoQ
3+O0dnr1Quu6BJkTUfwbRrxmbG8Dyux2oB+4po7UIItFgpcg/mBzUDuGPjIGrFu/VxzL2q7O+Tec
4RG5N5jy0WzLwvmlykMm/m1Tu6w+UeGkKbYoEDUvKsGZOYAKIbctq2tojKOv2/9pgr85a2jBaNJU
vURbdKC+hZ8qNcfWlUmDH8uNqua6ylaGhAwNbqM1vx1x0WXbnX1fGaywb2Lmd2/ZO2P/emMC3ewB
TNMgo+4e5sBmtobDHdHW5SqTRBukJtsfjyGMGOIpZJ5L9dq7kxa6ZE/qS+/peJ6kEeHAiB140L9G
Usvy6MwkZXyi7NXyInthcfjMe1MpIY/68j3ZXRx10DWgoAI9SC9G37d97X6p9PyFWN26mXpzFqh0
Asc45pfIdwnqRXVhhUMh1gwf0knTQP2v4uEYE8O15rj4DBehMdRjRjv8kEGbhbws7WbyA5Gtf3fv
QegF4BinGq3j25lOICl4x7N+zbMscF3n1aZ5YH+uyGlKJiYpB0L+VYNVvVUV+Hn6BSPi1y7teMBo
lrufJTeHmOEqcEkzk34dYP4qTdGOdQeZDclZ/4G2Wg9Lxa/h9UmNWNw+IgRJCU00fPGHe+VhD/5O
QMI82FMQ7GfIyvE3oKO/u+uR+IlNQjOlUuv9ehT4f3VsrufHZstBD6/yr7F+tUFG6JV6yCz0iGCu
Bx/vRRiercfD5KBDDHd5VWwcRDBdosNMSmUz0TFoDoqGo7O6Ib2L6UjbUKdXecgI1Nw2754Joe9T
JuZknEK4C8vnwqxLTBBQ4bLPLScblAlFokDmRrbO4bbT3zIeuCANc/BlIC2nwSWxWLfyVFJHAigX
S4l2MTbygUrRwK8ovkUbRKKKRCwjta2T3w3H0REk+g+kac38mmqwoj2/AsXVkH2mHz9lUjrAyey1
hzS6rLrK4w6fc+1pdIbLVGsQNJ1wd52ZN2zpE+Hxdy9VSa87xWMFW+N1OapqzPsKE/hQhxv9jK0z
kkS2BTPy2oEVhohluzo0LQW3qGYk0gASP+cm7jITUTZfUZBAAIv94i+hv9peX16wYkP+HitGbbRC
u425db6gxqJOnhbtIMJM5Z+u/FwFNTAIj9jgnOlIDPWA2j/pEMtwrSpcWBtHdl3lMFyDo+tyEYiw
37HYqgF6UFp2qzhvLykVnMkftb6zIkIOi7JruI8jA3YA5fbjcMI0zGmh8MUB88nrhAaynARN1jma
P8n3luIqAB3fK5vVu2Ow3nwwEkykQOS6gX1RoicAHdBpb3ysv2RtBIHQY8+iFJLmGaXoOBIE4/Q8
SUTIdZYNfQjsJWRB5oSvpdn3OTykV2yXd+pcMYkb7mo8xgHAFTcuK7Jj2j3ggRtg25Io0nytE9cC
81UbFaZTjxAhMzynILjfIriUfmrGIi3fAouCFCs1SgqAC5E7sQtr1TNn9RfWPNQIEsY+BZutMTa0
0IBw+exJugaENWueoJykxrUo7TItx7d6IdU5vwM7RV8Jxv4jnbzN/RLdR+v74mLuEE0iOoARLSOl
ZmGRVf6SLg3q6us5TSgHBwxPsSErA4aTDgnrYuBe8TUMzevoYUp3k32sEIcwac7AhYkeM+ZkLllU
5wTEzPx/0PnoS02irahvDMBmuucdVGHarOtw8ZtdvO30+hL7U+0UWJKYItobiHTG/MPznDKZ/nSu
N0XZQcs5UZsL2MnBnJJ38e+rAVd268c7pD6VwQdnF0Ut2KWjuA2y7NpIaYov9MnrjUqCvmrVOkui
a+7MkEqkzFPZsypmjheNc+8FQbgy8WxgrzQyBo32NvjpNmZs/O3te1/Xi8M9RnChEjz1JFacujAR
N0n+ukeL8PZQLvdDC6n23np/lEkuJ9xCYFUyjvutz/YEKlIsMGbDvNE7q7OnktC2ykhsHPv+wuaU
UBPuohh3qWf8hxEj/xpbh7+usRxwQTh7byhNIVoIcsmam4oqR8zAYBCHG0JJbMQxoJtEIgm9EnlI
Z1R5sLlJudWIMsbikYhKzCK7iyfEA6B94aN5xzywph8NtUoihG21c1BC93VrzR6ljWc8tGnR4wAa
LjeRXQy2LfWN9G2wa+XBWn4BwvP3OVHWSxxmUakuM+gZ99TswoXy1jd7P34fbvxbf/0HKJkP2xNy
WLQ+FEcteYUSqhexdM1JVvk96RKMVFZn87+RsXkeVCWgnCgbqTJ7FY489NG8SBYxj5sGQaCd4w+t
WzDr1Im8dqDiBRc2bEZm79EuEnOOj5a6J6BYHu1axyKYEQFig21xFodoOGTY1pM3ekmd0CF4/brJ
z4IRcTbEo29H+/xUzPZdk9SX5uTnzIBSpazBwbDsMG9HHPgwgOexCAGkTjb3phUz66hMbYBGxHec
y/pRXfXsxqwoXqOx01zJoYPOPHSRFtPaOPKlmXFI88FPp4WsTuIfsDjv041B6uEldAmJjglYDGD+
TYCdvUczQkpI3D4Th9BnzYz/9yDTApjw5dJqvZB6mFeJDdTrDItPxdkvCPbYERyjQOHH6Npcaomj
BSYPzpyBF6zP0Ytb1r4Xo/OQFzBFZfIL4v9kB5wA2Ju8AKKebeN4mY3JwmY+WbCTLnoWuPIBuKla
PhS50Uhsoper8J6ztsgKnvyvBhbOmJvWl2jQI7SS8bVIYDhyb9NIWT37SuI3ekek6iJXul8WDgGn
Jc0xK9smQyRDggedo+1Yl03qNSri1cEC76HPDFYc9C2ju0RCWNHSFV+CdvGUZ7T/ci6DYRd8ydrZ
VSDPI+E0tU0j4tY88kctcieZkUq6ToOMsPFprsNV5py3UFmUfxAKMwik9skn0V4etG6DV5B0LMFK
/XBbKhYqTyUmUqmHHwgJkURtlAuhzj9fxj2hgRMpyQqndDrklIEZZ0rJX+BTClqefqUqcNPuT2cA
hkzQAz5iXBABSe6PPAyt74eCMdGbwo6DH4D7on6thj6hYjAZKJbXJOzsH0/nYl/DalYEPtIvMm4X
9bFiO5CzWnYwX1Lw1VeoiK9oZHPx/JQKgwofCs1Oxn/nC4/tBMaW/EvEZgdDvYZeO/7pfeDp/sg2
iQ7XEdZllVJoy6VYltQobPFdrD/lfBc47tnuB5ybl2jbouNU0enI+iMO/UMew5MjblFkRQ6YDBFM
ZBj93fDwNiQJkF453D5VusDDMXUXgVnRiAvWPHlZxsTRqoUqjm0HRZIalguCkj81818Djc7uh3Z3
IURfHhhHvsRvVZu8Ohu+WG6FRoNft4xr4fOTFNT+74oZV55B4dZhV15Py8MxpE8NHBGn5hgrMquM
n/0wxUNVx5suhHfFMDrFcpCkgfSd3LZl8LtvcE8/p26mIDqDi6LAEu41icVqck+ynsXbD1k/0maR
0t98AuosSpJbevv6WS4NY55onsv1yzKZ4fS2P3JgR4brLX59mXsW6DQmcOZxGEmaa9sjC7Ip8YT3
vrccVXnvIOozjQeprfPKfl0eNq30IxZ9KUfo8c49SPvVGDmfdjhhD8RcECCRX9FFrxqo12LzJ7cQ
M0UxqNkvEXJat9gdoX8d84DRez1t6aPFvdbKb2tGvajiZg8SamsE9r5CbPFhjitq/41I2hIJF8PZ
m54r9jrywTF0EYpCmE0pmS49a3pUbCJg8TJpHGVADvW8JzQGdANgtbD/eyk6LXQE/RYx3ROJfjBR
Nvw106+ZNI0JihB7mleUhJrXc3uaMFd652iqj76IXa/937F6pi5UKthe3eNq+caomaKUr0//outi
cCZabQenQNmEb8AHh6zwUus0IqznpeVhzFEzv3+Dn1cMSslULioF+laSfF2ORZCLPyM3l7IBTsfL
XgfEbuC+GUjXldAaoXOjo4Uw2dJ23tTwSIjHpUzjgZ5CYD/ki1CN29j+VtY6lpshrI6VG8moNoqF
hxipHQNB3c51V/a1fW9+YVJYgjjQHBZCcVTaNcEW1OQYKuDrfPCAeDjqDRrl8Yj8OUN0OGu3187M
1XLgMfJ+UccjkIud8QZfFZnyr72no9UNr1dza3VZK+qUVY4RrBtGxJQI2L12+o/BirGxMpeWPprs
W9ed2empIIrt4sudzip7XtMNz19Uk5jxCdXoyPx3Ltd99KZPD7FyooneGFAHKBJhLs3A/tH3WuvH
3Mm1tKFZnWn1A9VZUZAciXL6qX9ifG3lJAcZi+pnz4JZXV04xbiASpWtj7eUkOEbOkUkwEN9jiWm
0zP03/DLk72XKYPZVt39CWTTOsxp2C9RWMdfbz+bUMZ0nzppiPeCPmlqHG0AhhLvE7L2xAQrI6ko
ge+RheadelnjRkdin7U85tMiuhRMy59RW/MG/4Hbulc9+hk1ONKY5UpuONCWPxbtwAPRZPmNQf6h
6SZQzXj9+zHuZNReG/egSOOerv8SWIxTHG0IzA9K1zxrgNiXRAeunl7Wjw2LmZmBk3rW32kMgvB3
3/mp1r4tEO+pDM2ptsL6uWoGChhsCX1p41I9WEAHU3HE15//o23owVJ72b0fgXlq5TCg613fMQff
La+e+qIjMOSHosaLRsbi6703/F1fkA2Kbg2vAxJfzqZbO3LcHGJgRM8oZPgivWGRV38VleR6Lf4I
XOUmPmNwVAR9p4rrP+9b2r8nBtU5ddjqAn9YzyhPZoJWyXMj+ZfkQ6crxeR4NPVP4LLUngATTtaK
IMCj+IE4q+9Ta36Nzvb3CgzJfi+GYMvY6PHrl12VQW0D9ar/jMCyGP/vWc5D/nyEYGMcSoyVsTGk
YAqB6KLMc7T/kulX6DZgPQNDZknSpiWKrdhXiw67TX/bgdB05AhN7pSLW+R5IrCQmwkQL1DkxZYQ
c9QzprpHFzBsoY/xnD+lguxKJ5x3jZvbBQ0ncinacm8KSoq3n3CV2wm8uH4VXdkzHMGiKu/h+68z
9P3b4BWmLZj0fGKmon9A2vzo89iqTRwtPTrHoksaqB87uzLv6/lSA8DLVW8CKjieWMckxfxTPBxO
iXScoC3oHkyMkV+w8Z041JwuyXXrr5JPSlt3f/O/zJ9toFAWUMdFsm7PdQ/TNU+8uvOIpa7Yi7Fi
e6sw7s0sxaxfAVOW2foFk6sKPdE4elGg8o+pQVKf5oSD8Leg+bp8i5lME1jYx21v2stHdGRU8gX8
V9nw+0baFOGlh5US77E1M3QVneuXOfh7vWZpHYl8iu6PBWSdCbUk4/J0HwNfQvTJUclr8FiPTAnP
nYS+ATXicka79FlqJHwvoJBqeRbXbt/pQevq4Dv/bvO48Kxqth3v/Msicn7jeDBWKRYpsQjCYcR4
jHp801H+G//7FyvO8YjOYheHqpoJQKhDHbB105XCMdxYZFlySt//dHVxsppWrFrh472JTYXVJGeh
FwLTk05dKiJmHZsYH2aEEpNuNvYP37PhtGccS8xUG2IHRUk1tf9MX9t4PVbyse5rhSdk8sDpmn9t
ROvdmWVdlk7qztHm2UkyYUvIpVgEEstx9bBk7sjIojizN5dr80UYf60eKlkxJY+0pZ3kW5rC8a4f
JRcCzMSGv3QXfEG/RvVcAnu0mjGiYPpogCDaNB1nkj/EF1iDLYcIrbmq/EAOD8GihdZMNqRk021X
lgunfZT1Q7pPpJgI1u4WPpqFgUrRfHvUt4R+OATVs+ySsmbW0Puhz25ryvSIf9sySu3yqkMk5ovP
Y4MlRPei0y4taX4e9ZWZNHJND8vUgy+XTPiBnrBVwFrrO/q5Cjhvgx8ndZjOKKO3sMn4+Mv4PxAg
F+FlIj+yHEfjmsmI2EjBv6CY+sZnCnBu6fkHJklwqRSdOvsH+zwWeCY2REWVyU6RuDXc+b/ozVgk
A316XOHHPEVQ0fiNwlInKx3IbgQoqVfDWGhRgTnliYl/fJ2RA7fx3tUC4xudVzlul/tbFZxI/R1t
Y7I0ikDrth2VEmrQY95UqgZp9/p3Cnp2STG/D6LQcQDjC1vFfxLIVMioCtkedHAuh4rQyTecnpjG
wzMS58P2grkK+tJ8gE6e03nBOT98zc0ocxAFqcre0fLwPXV0L7HK06Ax1V9+N8Eb8C5IcgPXBx4D
gQlirrfyBCO73QY+4tZR5ysWjTnN78my0ZZaNe8mvMJui9h3xyD0hreYFnzQEHcu/AgDcJ3g8RMa
0Gi87nNggFL5GOyfAp6jwVWaQCyhz/A5YGkyjLGc/GagVDB8jnh0nYrRffuLwDuQmQ75nrZGrzQM
Hnc1bfE2ygFjvKspZcjdgfpXHSFdt1Fbm3PK9S1jiM/IWW235nK7TtpijkEqpAU4G5Ug1Ib/mE3t
HY1Xhvl/CHAxctFQilEGYQPmyaIpUq1dmfOZDrVr/SEw6pZXBaLm8qy7JKelyon3kNaRlAisxOfY
dHJI6RmkiPTaB7+6i68hJjTaVSshN/S7Clzcl1ix+3dFGNpEVMXhff1k1ZN37BzzPlCOvZ8QrP1p
wf6hXTy6i6qcfOIyTBGdBszPbjgHvmpB30zb5erqR4LHi0YyINAbxmrIN+FoD0kGMdS2IDJ+P5iz
3pJ7CdS4zJGI6d7yHapi9KqS+mBgyM4VIo8hVOWVXf/DgLzmE4BKZKTiFhMXkBAXcNMsAepl0xIJ
rvB8GbuOZyd2a9gd8QkvbYQ77S2rotSOmRBVx5jbEom5UgmpjyTmPzC/s22Ywl43IoiAyr6g9X5J
UaFNB9jITVS+XJ4YjfEQLXjS5CvPc0X/FcOnlclcxQa0F2l6sHMac9cHVUtuYEOfX1BZCM/jQMEa
+BWtrQ/EsSDWZ1Q4/GMJwgGOAGhxz9OOKE7qVNU6FBF7fm7ShgdfpHtfrNUD8MEDJ3+LN74GSl2p
xp3R0+4fEuKcTmWWdELJKVYjbRp0yDZ58FbriYQpWdd54MgmIvBMML52AQKf0TVIr8d0AmCR6E05
pOrZQ9u9KRLNVe0OB7vMcDusGbuIF5yZHpbn5oBur8X5TnbvtGvX1INz1TONmBHMIJS1Jc1LxoNV
4vSBg9SJg519Kt22B/8G1jS6ymh+Qc0E4ERqXIy3c8n7M4+Kw0jm/rG8CwxigHj4+hLbrkxccCi0
EALhme6vzpSmsU3VguTfyx5PiQAqquCnXHOwzD1qxVK9iuAtE3BDgsiuQVMbihNTduTu9C7nIaBS
N+qK2JgUNY2iCktloW4aGbUxidlsg/+T5FewJ5zyikqc63vdqmyx7j9Mjb8EidoGVvxwmbVyEmD0
q5/0KeBpj2ABWcPblnsMuVI8jHVf2fg6PEN5/M9lG7dlYdNK50UNq2beKLEUzfmuyhKKsVRWKWdz
/ighWmIumqNoqSNy05Lc1T0HkH6LJ3P0GwtKF5aR5RFY5RvdwW1rFvqZimXrHaYum48BTWjLP0N5
uODOV8pAJp5yVU9rfzl9RrjeSf5O0Ussu6ZPmyWw8Q2YvOmo82CiolhI9sh/sFTvumV5H4cS0sWN
g4vMo+WH8mC2fvgkF156RQlLytgmYnNIz9UHY4Y1lLj1S5vI2HAnFg274ATHVHQgjl0/Z290Lx+X
wlvAWVRMJ5H8Be5osFWi/SCNV3IXIIdfCiqs/vX53AJV7qTZC3Am0NTTm0ctfYH4V/iYEKSU6DO9
cyvLgmxls5cII6kP7bXiJVInjyJ8HtAEyLO8wE7fEMKCZOoI6FBEokgUvDcNiXSdrnUtWCr4lpMh
dw1D8vVL6gPJMC47R+HyTjhQDptevcQQvkOzzQSCSk6oVpCE7DmLTBJWmXx+kNW6mZzKE9YW/cWC
Zv56qlatIsDwIE0PSVl7A3ThCFUxzM1bHEFzyRgsdLpVZEMZH1g/UXjaGF3hkqEcO69St3yCjeWn
IAWw3VdV5W1wB427ksoQHHspDkdsL5ocfsdYyFvUPi1LHBUnCG6z5aiwWZG6X1SAk+/jvIy0reIV
/T40AwYiqra90UfNmO7gj3YUqTPQkgtw8G6jPGBrt4rS8lp+HWVrvPE/FOLA2/ghD3u564+lDSL3
h6YqGQsfDv+xKR23+C0ofuNoUoqXqu7LIsVtoMt0GeiSqPMHRUadGUBi4ckc16EKgTFXerFn0G+Z
iWrOd82Mc9V14yZv4K+GuXLLkqQktyj+5iuEStGsckOe49TUr8DDJW+lVXcEpjyJUrYTC2CgLYsD
DcDc7+yXOJ87eSxLkokYRlB/8blxDA3D/z4NkwxnQqnBitH6OhSO5r6ebgEoVGvSnJ8gfe0N63Lf
AYnsKzcr9d577BX7KbvQ383ApJegNj0EajQd3uDxh8sk4UlVcVb6pub+EJ4+jGI92eQ7IU+BWcci
M1vcXAXPUpcFYRnr+a++ClXvpeL27J02Y4GbgIprFCNceBZ+mVkezgfEP8u8uxzQepn23Nmq5c+M
qblJdZf+RL/zW1BnnaJgn/+slQ0e4xCi/rOKkt+sGQSix26tnCd8OHrpEu8IHQRPSwbHV0rSbUYM
KhwjKu0JizVibakLtA83bYLyVAPiAwthiOSDTq+oWy6IEkqy8V3/WqYJ1senQdtfIY3pvZzKPRy7
puvX3tPxatFRThTMVKICz+3qGx8mflrGsdYssL8hsJLGQdKnctVjgokkliNUmkODlmL+ythOKRVK
fxr88mXqi8OQ71z3evH0LCivZZ3TaxysS6ndBafr0iUR5exNltlw3Mld0h7k3T+cuSBzOMru4v40
r/oKh6EIvdkq+OXA7jkttkQodWYEDpoAXHgTzeItJSNo7uLMytehY0jzilp9X8+BpLUnrqD0ihn5
b5Y9wV9njmHCSIenMbAslkG3UB+ZdGIVVcKrwYYfeNk0pMQhwMmahHVqZsfvzWNnlAemow7TmfZi
NcRaHbm9ez4+LSUoIoKdzWZD/CYaULTVPIddx5e0NRECip/9NjpSKtW7slvo+NGHEHJoZ0n4QuGp
F5YbYacJevHz9Fe8LyqjQq5tMX8zdVh2+Z7bIycJjzJiMs2fOFpBvN8tiS6IucK9uo+T5kDUTAKJ
zgfpV6PyRDLvbn1yipaCtq+Bzx18pqqK7WBr+ZBBYr4+4VxQhAaXO90gdXd5YbjXpO2ZMsS8Pjwt
a8aGeNG/aN5sPWB8c2uxQtzaBxnFkjp/CzuKykYRSCmCZamUU0gcOYGwAV0ec+gHVZyWnrSZaDbh
VyamNaErZPBBemj+RhAC09nDzEULSFB90pOjSCdfhuNEuLr7qpdE+RjyObqntStPSPrUjTBCseVv
l1tA76WFL7QzNYP5EIlj4zyXEvl+gBEJ5kRxyGOBu8mywQ3leQuVKP7bp7Q0/Er/AmPLSWvavfhi
onxvUbbVtqurx+RizLKwUbrIxEm0KVkJdIY0MzaaXXCeReZ909j8wb5bOw0oToI9xboB9BIkrVns
nY7qaYW2dcSGg8wMxieTAZntiG9yJZfV9VHaEGeA6E4KJWTcd2PibZi7FBLQcq2UgC/H45wzZEAX
M1cz0TiyI74QaSgkoMqlfucDBz0cVtAQ5D9vcrEUvCoP2tRPtA+RsEN1bn3zS3nSdcyfjww/1Nvk
+OvAIslVaAnsZVWkMWkTi8AIwH3mNktG6dRiMuedBM31KXGFjPMrXjWjufWugYiJk1hbuIEsRBUB
2qjetAwrDjymhUEyUcj//PfEkrpnXh6wWMMhDTWy7sFuejZJUl+RPjRddlGVdDx3lSizrAv4YaIw
Q9bMWN5FP/DdatSOu5EhsNd0yBJqwWFRwQisXDWG59v8mmG+flkbL+MI15vqb5tZokWutx2QMTLe
FEQ0VueHAnjTev8UqbQY67uyzDux3IbAqOuYp5ocMcjI6Uw02pyNGndIwyyS6ir/QT/vZmPolB90
3lq5ZN8bagEGkYVjsdLOK8h+5Lf5LRk9PvygayvpDR4lLd5g/De9tmWjWnUCcB8r/X9gmdy9rM+f
VS2YIfLWQrEZ3d8RpH+vWgVKnH1lXZdijpFQgZkp/DcEPXlqyMgQJH6M9ZkXbKIl/+0ePYlZlmbD
bKJirLjeQEzul2HPKmx9OYacml8B5w9yDZ0dAUzF7Gz1X+nuD+9DHB7FYtFlDLJAnxkg9EwB/5AW
Ek1kan+4t/XvVdEJ71wLF/UPjxmktNmkJy4JgGPSKlomxSN3PDM7JT9n/c2DSCfGxDWR1ADvhoWl
Rfya5Hr9mHY7KKOXWkz3AoXbLzDkfhzW1NdqsJzIophparwUoI5s8+LTh+vvYgDTz0VT0wuc/DAD
XlkRq4Rhy+A3RgMgOYyYJsbL2RAsJH7E2ozk4Kg50EH52shT1DW3ryCQqwNpWKy+OWnjTGAU4mXp
E5S6x5RTMrJPL1173Z1/MXC5Y8kDldl4nT6NTYtX3L/fMWzOdFY+MF9dLzN40KSxVYP99xg05DSu
AgN8A8eMBBJtLJsh11SUp8MA30420HctRK6RqOwYmimGnM+gm2xxET4ISe8KHtnCo6Hq0G4WIpv+
wXpuXjA16kdX+iJSJBzr3D9W8cptOvtq34e+FsHf0wQYn/COUpuoChL51XXeN1+Qb2M2PIis0YZW
rm+maFLPe4PCUmcDtYa05DTNEROvVDhPwWohOl0etHOZEibMCbdc6manoipiCzsSfgABgFz8frcY
QAjPXsObZrmrkgJGgDx15845F8Wq5jpNeBg2zC8xlAXQoGz9FQP3q0vi/fAsrmSfXVidHHdA1eBZ
cswD++Mj0qHQFtkrGmV4ouCh+re0T2MqrKdhSayg9ve0du2fMRT8mZYi1jvyJ+EdxkL0YX42xhoE
MQy4S3fbccpUSlLxZ3lasVTt1l8qnKhlk8VJVMxkc01JXkMi/GPw4bzf5JyBhl1Dx4ukYQpCruoD
eRobC/qGxFVYgvAV+z9vt1Hupqw9tlxLHi4t73DKcJpIa3bU4WlQeANMgh66vjUOs34FmbWXCs3Q
2cxt4lEBn8zb0X3IazJdBBmUBqADEeG8bIJq0/U6UIBs4OO2ThCYVUy7VttI11SknGTal2wREUni
W47AFY6ucJy1t8f8YJ5O+ttoDAbRZXFwQPaYv+vnqC+sVZYIeSWn6rveMZ1uBGm3T8LllhWJY0Gs
ojI5BL5ijN9tytpNMxtGRutszxpnXdORCf+4jCwV83lGRoXxzYUJU4sZFrKHS7N7fTThP6R80Gri
KmDT4bHnHB7lirXl+n5WR95LypFMydMSDtMhsP7ADhYjzWctBtcFMx6HKZuSCvAfwg0j5asCYrXH
eF52s/IY5bZ/OQgTb1WwvnLY7z8P+uzy7mWCyimpEMC0tA7uivV1Nurl7dQVEKGsbuT0GICGWOyu
iXoIyCCDixXpVTmjX0+dbgokfrkGy/G1DAi6as/yvQDyEIyMegHNz/R3tFHIF5IEq7NMgXQSg4pV
2t/pbk3TCzfoAysk9I1nvEqu1sTfSlBFA7r9h0wUh+w8/Nhop/krcGyWoTkzBAhdvv1uGUQy1PXD
WZHuT0G2YOmmwpKuKUw4hNqIu+OpnCMxyb1bE8cVLNjNvWT0EY2EBPjOhF77VU9p6fAWar5bYQgz
4IyGPqPXPGi/frW7orN817EpKz0VZcZjabANJvsVhRgUImUZDAlmXrI9Ga+tbkwUwv9B/7vZY6J0
95SO0RQXxcorh060x3vTfvnyS90GxUqvqIJCKRU0Fobx3XT+f/ZEOKw2ZcPn7ceT/dBEqHuEzky3
uP02ZWPkBEJSNLLD2Hmzr0OOQRkrf0zzQCStPQ10Urd4GDLODvLnjl1EuiriUhNUnO9oQQgT3j+l
AkU8Wq8BbAyyXccRwy+amz5P4O3hK45vii4CXHIqxFQDZeJumCxO5SzCIiNVmkkeWorVAXzzSTOI
avJOIVs/FXpwhzItKwekn+mepJO6xL5LmFovIBT2AcNqSyZ50W1wvC4KfzYoeJ5QYr9brwwrh6P8
TF4YXc9EIOkWMpD0jRZ0+eaNXkGtTQ1gEF8X3EKaGyqj2iuQWjYDLaknv+trPQmchL/iyZBue6nq
yT6zmKAWmH1el1oqfi55luu5WfjUQ2RQZFTkITsjmn94PInMMUZrI3S+bQKaqE1Z1AhAX2xhOEvy
GZggts2Mo7C0N5gxif4bChhz5nHpfzK2wTBJLVrp7TTwkFgv9gYYOfizA0PSGV7icwGcNAA1bOen
eLRmWx9oT2G0gT9Q3OMvspCu06xohZevpOVcp/clYoL3uVu8Flo2OIovJLD76wxCD19tREq1Hdc6
4elxCcW7SvEyLUs6YqVanSp3CFS1lRNXtkfs98oOQR2xVCzvhVEdzqVr6R/1si2erMtVI6VmOiRr
vIPYxw35zYExem1Hu6+EbPWucGVBmbo0UE/83kTljw/jxRw8Nfm3Po+6PhswzHHw5wqZvbjBrc3g
gH+crFbQqXVAcakHOcfx4WG9nkCUe4287WG+e+t8n8hSxsaVnn+d5fLDwDic8rVwtDINiTbd7F2P
tYuY7XRlI7G2SigkDkGzmj9J97SviwkoQOD5PKdHy1cI5LIM1ceCN8X3nds2ga0qMx1ksyitO9hq
c1zrAJHhXEaKMG55dOWMM/XZ1sFhmJZ10arx/SXASfc+rHXx2IRs1kceNu8SduBcYm/AG9CBmCYO
osb50jiMd1b6/2uXlUY8tBKwo+KHftTBgjAkQ7jIJA0SItsZsF8mrQ3gpaiq95qYpkpug8oFNa73
tj3dCgm6+ZZb6O/KTMfzyKRFec3iiLtguAitMszGs9hxzHGMp4f1pJGCCbRqKZxxFKcqhpInjmXr
CERDxgzU7teBuK3dj3xyRZ1RmJKHtyAHZR4F8a9K+41vjLILcZ6aFIkJa3/fBLdLQqPmMz3CHFlX
z8IM3EqUPGLQ3ve2bq1S0cVNqXN863DukZqxhZoFFvJdIrSjxHQQmoXiV5EYC6r6Hzv+0ngl/nDi
4lB3qBKBN6Idw6v2dZ9UaQifz86ItsvF7AkF3vnbU0cwuHo05lvA2IH8nQUwaVK7WY3wfilbdZEB
/ZBIb7joMpUi9Nfs3SrgYYKrjEHVkUgdohlYyCIqWOmaaK55uBMEOYgnsDSha8yhoiHo5sR6Y4+W
w/Nd7RBqPfrh5B00wqc7YrxnNTcmviFNiti/GKDy2ESLyDBPezXl5kVXEXaMoVCvMnjNsXO5QFjU
0RUWNRAVV9GMJeQW4rbClnvEcwegm98H78QBUejxeesVeBXMFwHB0mD+iuLHX8msFsO5gn031D5/
K165hAiYT8HU47n1v5HtSvug+Op9QC5RIa0GJrQjOtuhxhGeLGVWm/BKJYup/zYgnv9X5boNcR+p
dQhRcsS80Ehns4mqdQnAaSKOsRHZNICnTuEyFwu/ByWNS9nqcgyiI6Io+oHRy7WdU6uzY+HYPRbI
7czbUMfEG0F+/cXXSetiu1Lkw0TDGZ89dr8ABdmYmfuT7T2kBnff8ol8aQUEG7/yiUuTLa6pIrai
XqD2+PP0+bnnebQ385pkDIKtnlZXMyRI/PT2IayfYzs1PihlzRkdZfPAbHDy50KSUurI8RnXJkDH
bMCskEcT6Yqcike5uelIDTl1aOPZRE/mcIaNdJWJGsO98RQ4RxWQQIdYMC/RKQlXVO8eEBGv5JJ1
zuwm0x7gCU1c887CiiqVU3+4EsTzFYmrhZk7ifuipva/gFIiYYZ+PUlh5G0wE7DKzUjtvtUETm5l
p/j2+ME3Q0ixGBJe+Evapb40yX7OTkBjGpmGRKdHtbPTxlmaDhZ+tEL46O6rYyUJ8EhadJM+mfWx
jEaUVWkK4c1be65T0q0rXU8XwLMnT0hg6hPkhI59AfybbISEMB7JahSlALqZZuv3P/bJAYbv0z98
qo5rtvff7jYObwYQQ1dECpvGH3T8aWg6zdoB5bGdp1S0wuTXbx3mzqddAvjoz4WM7AIAZnQX03ml
Qc7DJEVV+/+lAy5IeGVQYhFOMt5ujG6Nl2oMaQpJTuug+JPXNX+MSzBn/mT7vomXMesFvKGmcJri
jGw78t+PhhFJZaITiLggfs4PYI+Utzr8FK/lCkxBs2dVfgMk/3tGgyZVqfdrW9eS32HPZtqa/NW0
Vtw/JfDNBdoQnaIetuwD3MKRgXRFoMwSrj8sY/05bax1zS5G4uT0/1diLRKJF5ACARoHM13jfTKT
5grRYu80qGZlte43ai/W6i2SVo5KBSucHXr6xbVKbcLlOUeDDjaGiu0V3kZv7Dq4B8dL/5h4KS7S
S9SYrkR0kk4gxI5AAz46F+p8eUYXtXRzqN1gOlEn9v2R7AVPoIYbZ7hONirEY6AW17gCMdJT9X3t
H1R/ot/8PVfSVPZ8/GNVTwDKivKdJIgiil65XjEzD0kPIlEQyhr7lKELw4i2/O3/EeeeOWLb1q5r
dRnCCE6kJN+vritI9sKzXz/2mHhTc9BJNw5qNb6S8EtE+symp1N+Mk03PY8fUzanUBPCJu2M4i3V
SSMgSUl5bg51iXemkwkOElljRd2JJEYBmolya9xaVMKflA3grgXHEVB5MV8bZDVet0Y+G3AKImAR
zSEpQDfwrn2ipmIWKg2hOff0IIZHyw+AQydto72gx5DmYaS3/S7ZldI/7v210VghdbeH+NTmv8VZ
MdHsZX1It19MiLVPtoMqF8Sk2lZVcMLpTROQZccJVyV28mcGAdlirFSaidamFe3C6OLPcqfYRvz1
FgSLoldIRi3YCAviDUjTTmBfKwZtVizgk7zomhWsEOeXpEZpFAhypbgumw+X/D5989SsqSBnNUdb
oQisrE8bE04dv99Os+jMf3xK6aW7bgY1VF0Xsr7xWIlFRu7sXIO0KpuQihc7AQTfWRMyK4NgszNd
lTvO9sGAVXzXnTqNdNwXGANtBBR47Akfyeoa+RJ/Zu+ZHvmmA5X/Pb73cLFkuobqDd5nIsilEw3e
k9GCJV1LRrYBW4a+dzbXLzGlsTyimI1waCIoBb2WpG8EBPAmZc8g1pvphOKxGbDX7ZCH3SUNYVjW
1tYzLSlxazQ9jInvbasnE2OVmGrj1HabvEtm326S7EW4oBE58kdXavyB5Pf8B0y8/QgI9DBqJ8D0
zGeM/oTGmpkIzpB6oCWUCNScl+ZEUiJ+GnzFMwvw891NeMk7MD9ap3AbzhNQFyrzRmQC+gQEYvPI
MNsN8UhaBT7MNuOnvU3HvPSzs3Ef9045zoM9Y3cZgsi4s9025xlweQFw1RZ2hckuIRyRR2ZQhL+8
lCF1R9TRWZ3JlNH1sd4oB8A6KdtCaZI5D9ZljRn5kgHxeZddnz7cfXuVqq8zLS/kIdjfKotmvzNb
+Oam9LvlnbhMxgElxv9gcCh3oGAPX1W4ZCtbTCKOwRzXtMajf7cxxRS1mjYQZotxmEt8Dx/XixdG
5RyUNjhKLDnN/QzhLckes7zxM6cYDHVGosJA9P+INkEwkEbJoyPZnZgHBdLn0aaO90kL4nnbdnRM
7A74W5nVigRKmEcKXatfmLAvc0Qty0TXW4e+SRzRRyg7YxU0nVya3lhgAccGRaGNeH6A/QNQnBia
GiMj2nEAZ/Vfc51ONiKJYP0i7qmYUcK+huULE+oRV/C8DDWZg1jhAQWPrM3KxMFA2cmkcoTdBg7T
2RzPnRIt8CofF6CwFa22ToDyBAjkbBBdxlOFqQnqy7rwRXXMHLMGWTO4NYDSkGt67crG2n/2UBRB
OqReGkc11e9LsJQT0tvZtkgq6xmko5IHp4dox7jUL7uyM5+ILxYotdLkql/AHjvuCRj0geuD8SeW
MaPJVyXUP1Uwuv42DZkzVlSnovBcqM2dnH2XTeg938XCpfD/MfXotehtlSee82DyBJqA/QsTPtGe
6MAim2hXF4pMjfkS9A7GS+lLJggZ5XCbfrZHQ8W93y+ol4Mxdckyp6IA5vADYlfjuxr5BvWoEliw
hUdMH3sQqRhPlGfGVbVAGigQMc9kYmsmAaX3HdW8gPND2j9JxBYqVkLTlzAPDMv62kHOhbMR4Kt5
F2qyfhPc/iZRPTUH+UFyJ8XlHDtSCc490RnaRqJAhLt/T0xEu72UyxFcYPua12eI2KuE9J66I+jy
9xDYcxakSxU85I0Bq5PhFRGCepFsHsXG3ede7Od+bCEI7KYaOXH83NQec3iJws2M7aqG0zmMhVTr
DYApm5OCQ8F/g0VWtIIrU1v3ZSl6o/cR4aOOcLSZ4rehCIm3MLhFYDzelYr2L0JuxEN0tv7iWKes
tTdSdRvhoxlCAu5rYpJku9zG2XsFzHhyTTrVyvPctIjQpsQw/L0ESZkVQ/84JVWJo0iWq+wpooeJ
GJXIxN6CIswcLK8+DnZ47hTQIGWpPEreBlViFXkH72EINC3vy1187bDnONomcY4lKOcDii187uPW
Fjv53IFVLwZPnLHijv9KxSZ5aalYY7uFEXwYttWABOo7dR/l2TxkMsCFBpJgZMbE96ar2MYoIbbC
XqMU7IADuSIIT5Ja3yvfQ7idvELNKwbUpvY4ljuyi+/jQAvpfiImkLdbu6g+sOUtAPgwTaH3Pzip
LW/f7jIP3BY4YOd11/KJORa5afgx+Noz9Hpc96jxUsoke86d2rdXru+FpP6/OsKFiCNFdysOk0ey
D0AWHuzT1nCwGedZwndypKf03BoyI2YJ2I9E23QsDUGPNLmtcKiwv8W53P7Z3UFSBRWqDEYDAB/Q
CH9dUZiNhqJhi/DjVhxX4mhCQbGySx1pb4/sLX5FbEi1xhfDY9Z40wrxEEDPBqpQL3dp2oOJC+WT
VtAWNLC7C+Dxql38rOyb0BBiBJqX36oe8ezO8pCbAk11Ekk7pEzhw4khQTroRCm/1w8bE/pCHrC+
LzugkdyK9qkAHrRw9FFyIeby6kc0zkE6CM/n6fEhTIcBsG4ik6Jd1iUwjgsNnHXAX3MYhW6HADo9
U7mQoxksX+LlNOjF7Mzir/JcfseEyu52W32E5nkm6tDWLDlCZQJyTIiw+PBWYYVnwP1zVPDZUyh8
S3k4KsUfBXpy7EWjVdQSX7VcogFbGD68gJM7OhZZbipBrVAdwoVJfjei0joebkxxQLBw+wsXrJ7M
jAdwfRYdLKlHknEQ3x5K1RvPKD9BZxkNM87ImUzYNYiWwNyUm+9ZaLL2KUaExxWk4o6SpbQQxEqs
4pNm/wsgCYysLx6q4fylapEYCKvVF6D0Oat7h2j3hkD8V8aZSHYz1KcQ9WIKwc5dQU41tcZwke0F
gk902T5OA0KxwIKbo32pouWxHwUbZervGTLkXUlqBOMxH9m7Q9v4lU6wZxVt7PboB61B89DvNXWH
/+KG8YS/nhfHyUuu68Hnx5OQbabsPcWkbeHyOupDluBzpyKCJEDN5zyPkZh+ahYDHFDXmWn3jVl0
aLamMPjliPdfehuUWaQqVbOmjveUsEgUbfcBuJoD40/1rzL/SudwaqcyZiavAF/UjdThI0FILGWe
ocNSMNwXPqfPOnJ2XkVS4K/JNWqD5RUEVJeldtze2jFG+/CfSr0410LvcWUR+xPnzLkUtKzModyH
kG3ZhVeElORlW56DnXLI6Y1UMAr7T6bfCmuFF4X3pf9WhuABIwr+jw90ETTaFN2v/XsbHamtqJRh
yhsDxlUTZ6lhmjckZ8qltanuNCVfhNDQ4rxcGsQFOCjyCZyEg1rC4SgkVRHHnrdl1fRaw4V6xHxv
icARWji/mJ0S8jGmxUFX8kdME8d4JONKlBPgbl7jneglinHi9EaGMi/cl49U0oY2+/WcDNS7QECX
Xx0HCJm/9dnw5R40FJfg0TyQCsuI82TbZ15DeenzQfumpYVGimMjBMkmjyvCUR5qIV4lrU4Emub9
j/7GogEeRpzjbNVlLEkul5Sop20kN1O2b+Ifd8aqbNFhx0p4qIgIbmf3Tq6qvAU8Ut9Z/1At8ecB
M+b9yrVC4tgNDqtSn+7go3YdBUfGK4rHXTmA2CvTA9fUXAoJVsTRTrqjqE/RWQbDGC75zV4FljQK
MONXM/kXXMmClOQ8jJKLU3gV4LPV33ardlKnQywcSx9QOC1E4NER00nYZlfxEb7NXCTd1Aj1A1mq
KhhmZP4w4Inali9O6FpaWB8yRoSo4PBkLyxNQNxGxJdbLPK4uYCPsowUU6e3SebuWowFBiRJ7cUw
TwoJq7Ik3cJvivs4+zzL7W7/zW3RqorJV6ZZN7UohK0hyoljJ70jdCfEknZ9XN8YI8sWwJJinPU2
rm0yQophxdOehuKiWf4taOflSqZtZFUbrXyDDyZKwl/x3jAkZhUj5WkAGm/wc9ACUJegCmR0lDJ5
gVxGvZTYeufyPMdme8Jy0gksjaYYH3IWE4kPcSQrhYpJ0kwXYhQZS5g/1s8cFe9/ATHgvzTjCe4B
MyqGRDgK/qpRBH0GZdkIsO8n0TYAhqenW21Pe3g7bH7b4EDv8h+lwj+VMhKavo9TUC5Tee8J5ejD
UUiuGvEdbBmaaQRdne0W9MseHgOveQAK1z/KKvzJLmoK6yZLgnTgtOsqFC6y69kAKiPu44j9qn0i
eOe8+dy5Foa8+etOrWCt8GVswCX5U8uT0HjJ6UZsJ+Nscae0GrOa8YLz3qDc6DDP6CAIG/YKRvOE
ESdh1vcF9b2b/qeIiB8AV7VmF9/Kd+3l/MtNvcGG96gz57Lqbyv7WvPUdc/Q5gxg5PcZLHm9YDqp
gsul2CfAJvu2eTdkBscWm5SEQ/vB/ke3B1s9WcoDympmnMpzm/MtfwSU4rDAE7xYxLUa2bow/XAf
oBIyc4EnfUo8vF05jcXkMyKg2KdShA8A1DbevnUjUdZVNgRcceKyyCP8jOcySWR9hqDdXkmqeNu9
lKzjlvQgYbfQ/J8sTCJJQSael2tGHV7FOu4ik6sLaCfoHbR0vB94q/hWENABRaMaXYu886yysWjm
8P07jzw3jwz8SigpZbm10Grp+SvLWCGUe5ux5my5RIKseUtDTqro9HLq3CldB+9Fl4N73MDS/fQK
k3utmpRrk3XWmb3sePzIkuhF6dnO6n6ajhswePL4jaUi3DxAh9fVRJyaCiUFjkoC1+bJE3+eW/h5
TUxa8M5WSozDlAmpedRJW6hydJPxmGlXLR62baF95f0ym7wTTuJSayz+O8hRNXHbWmwQZb56I5QT
xz0xD++KN/BIlEDPSksc6KAoDjTTJ5Sn2V9OmrrVbna2nL7N9uTC9l7CNZp4S8AcYBonmWr0xFPn
Y+NBbpnpcA4GeJKkDI0/gm4t2EUrrGw/RUzcovIkwWipkEcao95eqGJhlKrdisG0GU/Djdi+rPub
axEovJNRwvhOw4pvjSE1/xqyMQjjtvvW+MA0T1RaYhOnb4LA/PHDEneI7dGlhbhJModlaepDyyVC
9r5loihQrQDDHBs28cBHmsTiD6w4hNTdHHwKaDo3Y9jYuU+fufK5JyMNi4cW96onRJ1Fh3xyJ1Rq
IHL4YG9Er3BALTxfSgBmwfAf/KqVKnOOm5JDq+57rSGIOPXVf7trO1ceJMyj85OnCaJp8d//lU+s
KMPvoSte8eASHxoUPZqoMO8O5B4TaT97FR786a9toLkDjCXs2pSYyNxEfE3p+AWpPZio2lSr8Gyd
ub8T22yw/EIShdwczoJyLTlHP0DQ26zQDl/0iYct//dkyr5YquRWtQ50C6yV/8YQ+YggAuevK3jY
a3ij5fvfDtlJ+wGtiJeA/XeiYG/pi9lxaiWSCJVUp2GtOVfywe4uMIuHHh1/tVesO6Ah+tunR3U6
Q00pJUY1l3fjoQxWcDtQoxAipkJ4Ci558AHljagc3yLx61q9bX+A56PYBEf5vYbhp+f1KLmKWI2r
BBvG5Vc/+w67ciZYs3kLnmApfX90V1N3igxFRlUsscmVLtLzMj+JBNVcYl75EaCONinNKBnHWHbz
I5+eq2rXNg5hsJGKTnzb6K6UCP2OqZGRjSfMKmqCaV9QFjpDEU5nzAaMBHIxXpCgqZ5Hwh2YCNWT
Sq2XnZFzy8ly52fcTicbuhwNutEaabTmVGTR2/qPUJw1HhqH8QOD7TPYFLYwkL8uQXxtWEkJds0B
snf5pcNlaez52zuj3ooxMPV55ZyF44IET5Rlo8at9DKvFL7oAOFhntPyBgBEsuOg2z3Yq1Qy6xY8
eCuObch/HE2rarr8JiflW42LdMyFoQWIYcL/v93DIcLbBkX30HMlI01zKM+TxR1TvzU95aVow31n
U3a2lgPJMZPdwSIgM9i94+oePtb/J9HwtXcCkbmZsv5GVnzC29e7LgEtsZt8AXmQjTB9voRZbV0a
qzvT0SiEM+Bs+o4nbENi2UpR+HMtTK4gTHWmMGuGB3S1eftU2KE3ZeJl/lloBj1bPepWQBCU1xK4
348e13nonOvCdrTP2Os6GQtg/7xLrznWwZ6eMkzNMidHUvab+qn1+VrM/lT4VZ01ZJAOKqrb8R1Y
hJQPuoqUYU0cOLRC0c7Og888l7U3IbF+eyXCDlW45X0GDuyPUwkifMQAHaxOSyba33i4wqoJWIIH
i9MbvoHJSzTV1YD+/5pc4twovcEo9UpLDShD4u3YNDvziXLRFoN/gt1XF1sAB2rWnrQBUNU2P8gk
gGZbtox5VExiFaCPsxjZbZ24eNk/GZxNV6UGpmvenD/W0hUHs+NPvM5SqjwmNKA7ckRRl94vIBeg
aA5D5rbmG4KQ+I8pgIOnR56XHt7wyvi6Ut9/wBEYt7GcWFnUDHxMFNaMc0p5TYCbtfhYaD2O0019
MNLXGNsPpqJdkMhe7g5zG/HJfAPin6sxKCXuW78YTUNk+CgaBWc/3taEMqX9oQR+vfDwwEbcrNrg
zdeZGXf8C4guyTqXrumL7Qx6RVVu+KXqReNVu5rzmWA4KlhUSr8YwL/5JWnI2r6jtLu5bnku6I/5
BwI/s+h5jqPePN98gc9/lpxsuoMJNh/VPK/BldFDnEOM+xgzjVFWta4dNNQdWK1b1A9SdsX08A8L
qVfwggyaX0SIahwQvJcpbPR3lUD/qI3d/H3Gaj0YaXhDql06azdU4cQvxAiuJ1/z4NP9vy+AGQ1/
D1TMW1CKnCdwRBIVGyjo7OXzbrDOGpSlzkmvunWyKe8AUTmx28lCxmC2rAmHOiwusFSYyfNJ41ek
mhy+Q70u2w1GCMU6Cpq0YScnx/GNfaZrn2hbVbxVs413VRHsplQSTy/DLfFL7zC40thiu3WwAAY1
W7CBRliEZR9NZR9WPHRI7czoS9y69c7GLrPRgloA+GGB4nZmkG8fMz3HNW9ClLaB+J1dLq+y5gwc
ElG6vBkGiz+gYR7v165OtBVMIuYrtkFGJwyVJwp+WdJsJd1YyXSibxMMq7lQ49kS8SiQFtYFOnqg
LiMRM1pTl1mH/cYtYXKDjTTWMLkRc3O2FA2Loitgsu+11+SyXSRYkt/apg8cKWXfjMFgHAVPZylS
xjpmWdc2tep9WTELiiVrlnSzCFAVJY/xlu2i80cdcAHHUyMUJRLw0uYH9tiraA0M6DfVIjFZSkTW
4A7FQwdHjRCsTA67lI6qutCNcggDqxUlq5ftCSr3VRS9wZfh/uEbFrXpA926lTA4Eid/+tUs41Uw
accG/QQOILSsIKrkMVblA1ZV2Geye414Qxd6Bx528KuHta9at1b39yjeEChZLR17wAF8oNj24uiv
25by+C7kOIceSDis0RpcHVH1dg9+TCUP5Wpqty/pARux5EGmy/+wtTk4h9+dvuWdGMb32ql2Fbw7
9UmiVQZai+ZY+nim4TxIcwTBLBsbC/PaUHSh+bMwq6CMTNiOld+rKXCP5mEVFDSoy1E3/SEOMS/U
Q+QnWTLsa0dnNypLktaalx7gueMvrfBaUtA9CFHYl5LztrECAV4AFVF5SDOdg28JS7+ed1EH4Lvm
ihVIzApHsJnDtq4aTSedRe/GeoOJ1hKb+g3nBhMfP6yW4mi7EltG1gnKhvehUkedKfxsLT2j/cfN
QlBZsg7p8NGwg0CzABC72HP2APvbusaKLp1Wb3BW10r2nqaVubOWlLYUu0TlZe2lgL1i4iVM9GdV
K5Oc8uEW64j/y+5A0E6dcrQ4GQG3ZYB/J7ZWYLkwa8C4wqMxBuO9vy/i9iROJoxQvvghrf7Q4ag+
wNyNH1fd3C+r5XC4ohDukfbHsCvU1g/qDEJCXWGADQP92Sr7fjPXHDF5xtQ4+gYN2sbRqoeYT4Q6
01fsPXRcvf8Re9EUTB9A8kFx80QzXTRQPwAcqqSeZ11Hy0zMsbkzylE/ab9IF7oikOVVcyFixqSN
fwhn5NnF5nwNxTa3sR810BMfP3oIBSwjX6WI8vLiAyRvT12CvduDwhaqCXVK6/etqhvHbh/cJ6n9
joJTphjzBsKgSxgjJsIYiYzpv4lKKFjlyn79wykkOMDQoLfzdguv3LB1fRxIq6bzyF5Ufd0Gs+T0
rOBEYz7vLcWmXof53ue+zn8Cdf/HFojt0y1zwvlIXEsWNjqBCTtMV8sS5ttbEVWPtmLT9c2nm7Dx
Pd6hhi/1oIzn9bUERIZ5abqL+eAfnTWlycflW70sWEzgEtyTjES5sxAnNgrJM1vlMw5wW0w3FjnM
xop5T6L8D4wEQ3sU9sHMQ++IeKl/4oRlmPv1CVP481rGodJGwTx7Ek9XjJ1trioCl7UTO8nOG2Rk
XQEKswZL97GUdxbmIDZJLaBWJu7ySE1AunwSOghbBQZmP+4Rvlkp1xBtTjA32gBI4CJ+nrZ/L2Xj
KYSdeC4AGile0kcozfkILuE+Z+jsKJsoZcfG3OUhqnEsn4go7Vdmw/v//FC4/hapQIiLG4k7kWPX
h64aV+bLbwDg8GbnB2/QYJwthrWlX4mqyuyCTGh4sCEEKiAPxRLlj3r9K+Nt10kZA8gdENCfOcS4
hS7LbtgBzVRmd9l6/Af/yg7srmx01/8w6+et0xo67UeTYZsisUXh8i6kwj5r6xaLjxIovY+7ZiXk
CyQ1AVONppPnMcknO4YFW0kK0nvGULJhRkwThapS4WFOuzTkoY9x6yDmsEJQp+vLbZra9859mDNW
Dn45cg+44cXbDPDrU/hLr1KSLplpAqu242HghqVPmks/4sMhmL1rEqq5YdL91Chx/0GYJiUqj9KJ
mm74AlcHBiqmcbYOYMPR1aQZ1yxrrnPOBe3+leQR83C3X9G4guLzpD1szIuxIaqUXq0oFugsUB5M
Y8XvnP0aXSlxexU/Sn/hGsERdYcd0okeQDlvl0xMmjwZZixzAaV8j4GIAh4lwv1IQF80hbCI2kwu
VDgsKR6b9onoSc7rRTpwQnBrJ0e0CFnH7RcplMcQheqIexwyCRUntVWCj/yBVza897kUDrZHPMni
a8dzzEY8HdZowgfN3v/gq+hCpkxOqxz6czWJq7MpEzsVLzDu3LAOuy768wueYXlB416EDBINxlwH
vXrBZl7ucUfpAdj8EUvWq9vYYA9MjQEKmuNi6rgnbv76Xw7TnBGGQjBExCQ/y3BPDa2tLEK6NFkN
od6ABEg8UT27yrzn2W+Q3OeYjLEQbaEQdo4P8Gbi0eRp2DTBh5fzrPCrTtF4AMQGxjtP5bcnm9qc
VkzB0dr0YAxKye5ZlA5XqG+L1uxW5KE3xZjs+wxrJqJDELy4qYUkOnu50nFisnKu5mbM+eM1pQ/1
tFGQR1NxVP/Nk9uNostvVXWFzlWgM/AVbIG2saQJrMXXATjZ1j7FzBJoV0XWobRJgZKyF8YN4GPS
Cxj0Tfk6Ack3i+tUqad/moW+OvxaRV8MWMnr7QUDD0EuCPGCotgZobtUy31BwJ2RAoL50fr476wd
fNTNsCEK3zUruBtYDaCZ6rRElDEze31E8X2tp+VAchjHo9R5s2viJH/X1OpDPpkvq68npQlHwI+M
DlsR8fHOwJDLwMp7hhTrFSdW9OSXO3wK0Dy3x/JXMQzQMQrNcBF1XRVI/U0oJ1IVjdcTlSt0BO0R
KVOZs5EuQ6oPxciUCsYUAeW8pr2PSRVz7++lCJbUZcDqvJr0ZLqsjFSsrwzgmUfOTIq2r4qOmP1/
dzm5c2oAo98ab+H4n3jUtj58deW8CYiBzp1dtFC+WXA1+sOWLLaHy6iJmqWfVI9OdPNobWb/qRLu
0OSmxAWDjHe5Ck0gszAVJhC/HLa0wq9QCvHbno7vWq6S2e0THy3ARVasP5LUyUEXEBxFHbFgpm5i
vfZuZZMPNxGrVsN2DZ8nT6ZIw3y18XgHB9T+l8VfmFbs3AxXiULJhEi0+yAWqLmkLJ70Thcqf2GF
hfScPDkc4wtC0mhvjIW7oWL3bvZH/S0Y7iPgGnZ9RPKwCtnSGv2WfrDsBqRU2ORsdgPbGHb4HRgS
EAUaL8ek5MilaUSgqtG4Ud2Nj3lkPoCTz4Ff/mkp5sXXJ9B04E3jwFCvz5qn592g8wISX6t401rS
OLIeWaz4dPQ5YRD6vG5Xb1hDctT5k9hTSyk8duM+Ereokxjonyma7eDuFuOYcqidTOmBxu4KUu5W
2oSCxmNLqyWfI/Y144meyQIYtNBh129kYSLFs3aBwVpxaZ9k4Wq3heK4McjqWTcA23xtJodrGbyx
95Wk34aPnb+VjWHQz8JARMgBw+EngwqLtBQeBnr26kXHd681dpK9h1N8XwDh3LctdtPHKWtYamOI
+XDraRszF6ThHSNs9lAMoThLozPxSzx3PK8ifyKbognZLd4Vj1wQTfDKtFD3KP5LfUIGo+U6/bak
KbNf5/v8fDMdFBfSQgA4EwpRxdAoXWZzG048Iwu2fxkFVsVijO4QUJHnlmb5Ff0gZtSf/Ev6ADRf
j2lLL/0Q6NRWeZTDwQfr+fnVDzIM92vAB9+IEPMqSZpS8MOtNML0hjCDI8dByNgWm/fYrkA3GC6X
JSlTeMqmmYJeWNJgVyLpQ+Cjlph19gz/irmLlTfpVRhvodkcYw35oLgSaeeAXyzXyT06i5dZSZXz
x0bo/5qmO2epWbELqzH3vdaa9o0ImNjMjUtVQzhkrQsQMP9evEAjqQyY/NsegxsRIZ7cuxGAoAj2
lEday2gCkFjREt51O4K7p8nczn77U3PkugLqRZ3716dPHegJsuMqiJWc26ub0Zcn5T8K9eZkUKJr
zpHXs9rt100WQ+oPpPXRYNWxuju8omp1evrMsZtZqdhoHOXn/Bf+9Ja1Yj1oSRUqznBPZ0wVlLL3
b0yJs5XrUSD9Nxk98grZpMYa/aM/f1CfjGfVsf6iYlb74CwB74pNm8mrGzrIlftzY34SNrXdBXd8
OGDT6a7EuG/ew9Xv27LPrv/mFwTlvxnL7PbLiq/kwolciIKRCXihtu+VTByQo977thFBopFk9SQ4
gCdSD6EbgM3MRac7t3n/He5MF2VFwyBKEOa+BsHUHVHT9o4nmOknd1RALVepQWR8DvAtshlv1mBT
VqlOKpA6yEq/b7GLubKQABzaP8aF8rGMyt1UtNF1h3AtBDkeGFZMxcbhEhkrpYmuqrSOJqtwVGaY
bIfnxrrcs+noWs60N0OHApoLUfZ4MZ+u/u5cVXPjSOLeVRuxyM6b7f5HiTi0NqxZSO1TmkOfTeIA
74/9cxhvLyotooUYDMl6UuPSwMoZaF32GT2lB/dVzTqtqzRgbEcrWM++Fu7XjbSWwZz4+iL0A5Fr
JdR4TNxuLrVSpd6ggIFcHSCx5UEDIx1ahQi6cx3IR0/Pl15amlelH8ReiOa9zwFILMhx1Tpjgg7s
cS/DP6LsXEoCDym3+wAOyWslaMbE+jqlwoeTgA0MKrqjvq+s6N+mJ65A4dmkZLyfny/DFwUhfoPE
yUKJ8GLibwkmFQOJqRBPSMDylVN6Gs98lulzFrxAkesehvqC/qfWO6YhLLIbEg8pw2LP0GWijdNw
GSt5o+Zb04DBlEf76epOvUg7aijFtxIuyaUlRs+C0z6wA5EVwlRpEJxqy6RxLsDk6O6Bn36chXas
UFCGELQMgKG2dB4VwJBO5WBz/n4kC0Ok3P/zphb4j+FqmKtgNezUxtFJEnhUrlIe7IaR5ZnoNHtB
GzE80zoe0KmfCXLSRhqn1aU823Iy1gMd+aeKFXkLFoWkWytw4F29CdQLMMlvgmVh1Od2TJJR6q1C
6ZjzTIDm2d707AZhHZyBNFJF+BhuqmdhAKbIvdlwWKzCyoIW6gWAXlqLmf/C8VD8fEp4GbTlfgJD
nTFAqVmqd0hqeU9BVMtJwUj0Tw1ITPfq16dSlYEmVWMIz0PMSpJpGqh9It1E7BHLv/tKn41RE8IU
3xjLl7coH0GVfHoYW+hDjkuZ+kDa3JM+gIaHJtMBTLAFikYecznxa3kReH0pRMD7R7imKJ0hWITo
wERVup1Dq6F4dej2pbTeZcdpDtzGUq3k9vH1LCzUIvJjkxvLukQzdQuSZEHuNisiRX7vB1gYRJYf
BT3ua907fD+7UCKSQAsR0A76DmLnH7nDHI85OV6nsVaE/FI7Xb93Odx2dvQqfP47ToVAViVMy+K7
aOgxbwT6mswOgcyJ4YNud0Btw+SlrBH9FnG1k/eg79C4XdsxQmevLc23IWzJJJbqXi7vbLKK6dK3
dilxPTFrjuPIBhAXqvujpQqJJ0zIxhByUAXr+k9kM/6wZ7nwTrDMUCXy1JK59kgt+0/IDC3vxIG5
AFl6lHQeWAoq9A7r3kCHXTKITzjsGhTzrm1/kvSFdacYcHPaejEko1tizkWyaga/HikIxQMzyZBv
3nx/l2JvvP37IqOduZ6Q0tVB7itKEpTEmds9zLfeaxprk1jZumeKg1tUjdCSG1XR93ZywOpYEv9E
oUmUhhmunXC5uSWiAu08JmUqjXLAQAFs5XGlb6Qn3GnMErWxnD7IoUrJf4xPB4DDhp03QtLse/wq
I6WHxBN0+U9P+ILXC7p0M6zXO4zTF/aU7FjEFTTejALU6SXxRK9KllO0FvtEStHHTKpLd+WH2lNv
iXRFaWeAnQkM64+iTrLyVz+/wN9ebdn3cbpCnX4Cjpq9oosyCT48TrPePabzCamI57NOe/h/jiSb
ObHFL2LvWJhOdmH772GWjNQ4L1ZhbVTVl/VRihE7L3DLVjgMT9BJZOTt4OZoMpxPh3gQz4ZJQjkp
GHkPtPItLsYRgGxhDwu96Md/UD/Y2E5WrGFL7VAX9ojFSZvWjsb+QstOp4AhNWVHsn/JrWPJdlNb
puqDqWsY00eam7GncED9sYNb/VvjWqx2JRleBcCuQHYXyIXfiDmUX5VfMvRUPR6tWzmaubu0ZdXh
VLkKMEOGQ+0T8xrkPB8vnk31tkFzdafEhTJ41lmIdOAOGP2o1xYbt/LdPZmY3jwql6Btix1Szz5C
iVJjlDQUHPQeY3xxGCxrTwuHjiYh01dAp7xqX/JFGaHXvhi/CUr+VjlU7E4hlsQps099XB1Q9pvH
AaGNUPZ0vjC5rsZ86Y3PiwdE1aAP5dOvwn/03q8Q2ngyd0MiBxWBh/CHLyLhJ0LNGyTNasidgh94
g+HhIS4PnnhZhRL9eBmZMHuMDDbm0W1dwQ5E+F3GeP0fihF0pFLZ3AWM8W60cH6ywxxjQ815WiIb
IBRdUgJFP8zdSj2/T8qjSG+nsoTeidA7VeqlyGXgVKVyLGSM0XtXJYJ2ltgqPQWke9zYgc+HzUiF
GaJDeEaIx13ye4eBXOxGbYHNTkmGz0KdpzizOlx8PbZBg0ao6RAaSFNATdaf+Cw7o5GlQc2lPaBD
o2nfVkiJ7AocA2v4cn69BITnMfv1RqvCOas3ovm8kdsJpyzjByoXeELaJkc7+uj59trtooB/fAps
H1tpOU+zlTPJWD5oim6/9Rcrd3oJaCeF1ISW0I5AOZbkyLbE69PFVQ/lgsTlDKQ9Cg8WRgoBd6KG
6tOJBJROvY0RfCB7Dk0gm5ajcUnIaUyP905A2F/ivMs7MQ6Qm/yGBIlua38Zvl9JdD7ZsI4gx/nN
rpe82RJeF0CBUKx8qormychknZirO3lYxjLEEdCrSksKrFqXeyVl0TQY+sBnkXvfStlXTsrwdgAE
rVC6BbMJ0etA1faPS57bA1z9EFboMvwFuAFOksH70iF9B1dRidqT8u12U3/az9Hyl56/C9NiwUv/
tE+RiLumdftxrRhg5wK6rmPrs2212WJE3MkhF1JIMTWKTwkwkRae1YsNQ/mnQN68ALQb8iiawrLL
YOGYryUV8k9Ifd49MpE6ax+OCw2qAGqLMWoF/rZvHN9+OOdzcFL1sgI4TDi73xf0umLsJGhi/FXU
U1Oz/ua2hDw8Tq9hn6qdObFjbEmE5T+T41dZruD0Ya4GlqohkyfV+7r5+io99G7v/KzMbFAJCxV+
RzMrJ1m9Zzv3JGtJqVdMS+znRXTb+aIuC4HvJBXDlk6nMXSIF60aS7wG8gHgQPd5Pp9kJhPSxcN4
H7lqbzBlDy+N4FpSBgw4t2zL6eDCGeVx70r06oOHe+klRWIi80wCBdRLncYZeJp+nM4Xlh8oATAu
PzJJYQFasqqCV0TQNkF7wxCJc8BIacyb8A7a11FhlLMPRuUHbWahurGbpw/xg6IbBF33ZNy2POeE
4H6EcTsu2OHZy3iongOlokd1liPz/KBMy2VsxXV4S2l4x5j19bBXgW6o3foPrajpejfFeLQnb/Nr
0WhFKhbiFwrmYyRU1bo9BnAn/CkDCHdhYj1pGdFpZLU2iwOqyl+8el1RwkC2gqDwR9WHNhxKqZ8m
59q8kFQvlKEecpy4AvKrF/KKzF991jN0xOVx2hmSpa8EmMX2R/I8HxP1OhtVW5xTa9svi9TMfMQ7
ZMCSfKwhdPwUKIrmDgH6l+ny5rnwHG+/E94GBz7wSnUVuOmAT9FToJmP+YkJO7DCq0g7n9Z/FL8I
v+zRvG3kpFyyjus2Qz90WwnwQNP5eRs5crM7TvXJ5o5A7Y2VTWIPfEa/rNalxUZPt4IRPK9hd4Rp
9TpxHivo3Q30nSSWMF5mUFFeOIdyq/X6H6kQ65xVoK3008hv0ctK0pyyopLIv9cfX7bUj+krjHbq
NUfcOty01yk4k0hgYXtH/Ftg+xXc8SgmPj11SCAg0MHz7GsLLT7BM8OSAoJsUf48LpVCFMvM39y0
02j0TMr0Oiftq5ApBUBM3wKpM0aFjwbYZOc1epS3DG0RVoFpXDlJ6c/Y0eLGSpf7Cf8XrvO3ArJL
VN7oAuzvPL/9+2XZWYWV12+OTxteDf5dbgWdNvP1JD+X4hQ5yaCZh0wgz2GF8kUc2SCBcRWjk/Q7
TfEnxdcZhDCSVvYOZSHAT1ao1Tf1V1Pl44zZsZ/9+0gR8gKVbngNBpnvWUoo0XWyswzpcDsqGPoc
7NzURYAsiiq+XpC+2ehPuY9omjJrpJ1h6fn3KBjlTThR8bCxjLu1SjVr1hm104N9XaSOuP7LA9S9
O1UU7tVMMFKs4xJozFANIEaibYDx58jSOGgf3MsEG2VbSnAYX3srZaiI+tgXw4iv3OBr75qAJ22i
Asw2ycuxOiTMeMFa7hymO19ViGMV6gC0ZehmgSn81x66JmUdUtUlO23PzdywYOlGTIM7EtJBCCdt
a03wGdfDuY3WzqY4NzUGTL56CoU6INxIWttJHVHsDoll0d62pRmQvsEPw/2+jI1LAQtvbQKA5yoJ
hUHeeEjFkyRU3rYu1wti7Swp9G5md9qdd2OiJkuk2l8CeaXmV3WR/5CYuehJafVHAlPRUfLODNbs
jOE77N+VxPMHv4PWIJ9dnp1WuRgqeN3fAgUoNi2S/F5GB8HehKlvkVtLNpebBJTGgfmaF53gvb2G
HMHWSIfiT9Z7io2Of/D5hNeyNITt0m7kLFohWbJ64i/aepuJ41oJ3naBWKJasr1VcOlo7cgWbYX7
nqX2SKiNxGlTWuG+hqayFPZIyzyhjYPSoUsesyEJnKc+Seg2SSUF/u4cEKmNeB81c1SW/DGA8X76
RVGsHrtgHezJpUem/9GfUENCxFhPwLthOqj0MGtxam5vV1PEDGSGGu/U0fAniz0sHTyWdSbbSsn3
5Qlytfaxxylhtw27LHhaC8mYwMxH4S56lEfZ1ZKonFjkjh9G4b3NEhWKRkiIioOL0NnP/lnhqvBw
AgqwQ60STEiACd+GuoWKx2i5OSiNvojWOfM9zv111EkX7tTs3WH4vTXRMb+ImDnVpKpyP/LV8vZq
HIGFTv2Tc7EEAPP55lz7qZjnkIvLpaE1JNxO8r1R20OZaHt+7wf63sQRgv2/Hj26V77jsSGKVTph
x36gTE4FyA2TVOU+NSA4nH6h3ItDwwIEZWWZIjLQ+ncgblhtIUgQ3IpLquHBjBvfjIxA90i3UdUu
IVcGInhrJC9txvc/JX37ELcafhk2vkBPabRdjJ3GE03GLCD0OgJbPsRdZz2RCHzQ7kDFdr9BGTcq
em/RKenh/120qkABCan3oT63hGUa5uFOxLvTezmTuw0niz4axlvGlAKxjxPvK6WtRbg4sLiehea5
CcZdjUIelNZU1Kbe6wHbK1qIWbZiiWsFmBt9RnFeuYV00yBAc6wn9J9y3o1ub+10+NoUtsappIqP
bYa2Nl92SE25n4kdoDWXB88VBc8CxCAXEJ0dX66hJYybWGZfiMsWKJ9+88PPvuy+pMFttnprvkl1
zCAoAnpRYZFK4/XWQrcROP0haAzOEBijjHMOE6sIvVohDyVDsbuAKr7+/kIp0br2NNfoy8UCkXmj
eRLjg8CZZJqdrWHuuKQchiJDpctZR+c1CPeOljxi+rn/0KSuZWxgbOYIpC5GnScVo9scRDCpaE2S
P8+3lxmagSxaIImjCoKz+q66OGKLEonVPR9MBwOjRC+2+beQX3ENgV+sF7q2KWUXAzj4GB0XXAVp
YZ6j+2FWfHntjWY/g8wSuD9lFdPmaJ1wOV9wPtdH7TyTXs0WEbwPm35DsjXQ9XRn9sMQAdUZOs1/
e0Me/WgbQzCmPshpUJjkmOYHOtgp9XQ3uLPZiiJwpJ/WfPIbMV5R3/sQkDMIIjD2K3Mao7ItHbPC
jzJhOSwiNzSn/W0FNud+F8vGgVd+vd6gate+bE+2267sN/Xqz/3RwSWqdaNOlY0TMPsEGjuw/qTX
VOArKs5XBE5Y+5WWPFG0fmdUkBhdCGzAoXnS7WCfU38I3IZJoEl2E8QClC3uCJPe8F3zqZ3cYkNw
+rDQU1xlMyYBFPF1LKWVzSVHg4OpWDxXto7MJBnWePZFB4J6fC7MKa9f2cxPX41oXzJ1Umje44dw
iRW8XK20WSrZiVoIGbm3/jFT8VOnonW44BABoYMvyVv9L2SokSBEtlnm00Jug5riBHPABLI6VBxh
qkUfQ16ILZ1ly7VobMxP9KsXAJNVh5YgMr46OfFMgDaSUVctJ2tf5cGtyzOhs9K1Q0hqHH2GUNWg
GwfmwwO82pKvIyoQ7ozJL5tZSfC7JjpO/KdT53mZnGsuykcQbvGvjZVxaVpaUVj9v0lCkTvdZXV0
XRgylS1MJ8zMGxRdlLV7VfqbFiaBX6kPrNfp+4HfLWsa4NLfLxgRp0XCykxX9PP/HhEf3aS3Y8Ls
ykgFrMU2nV56SvaE7DnOZgejHNk4lA60jIvT2eG5ZmWywMW0kvCHhnW89+W1gu9WhtrOWMlXLzao
jf8PeoNmGsYxNy+I3ba3x8cAfUuortlHpswAqBP8N1SBUYqth3VhkGy1ox+0CASv0ofiCMELw0IT
CT7PGR29m2LR+6Wygwz9M+HdMSd7lJP11fwm6kakYWkquKuxLEen0zTjuRahd3E+Gv7VNNANnPfc
KY9GDtJEUb2EAWHJROkydB9Js3q3oDqardjQhZ5pMQLC7iOeMyVTf9bEcZkHyPOogvkyWRb8rRfS
HP8uocj0sKI2hghLNEJfxwt0h/uTidAa4J/W4KEimcw3FTL+tAc8+ZWkk0puIoXloUcykRxZ6BnC
918TFQkspzhcyj4R9Ar60Y9zmDTsWawHPiP4+OL5eGapMls1HLCip6M9CSTCyJLYPYWsRC+BUu8+
0sxzxpQEzMMAqIN+BeCxUdPaAO8bDWadiu98eqP0QSj7wwHhg8xGcnjAXmoqYmmwGUOuI3L1hjBb
leygieiHbShWsfqjyp8GPcrma7w0LNyS+eIzyJy+IKRRatN2C8Qw7uIyhRd6a8zfLKu45/22o8+j
3noDihr7cIWIUewzqxkcA7JsqUvnx8p9RYQ7kkb5Li0OxTa2PZoh2j3HTOWV2ZlBKXZLT/jTJmMe
OqPxgNG6KVlMnZH1LYqPQLSFY3kXSWfhdv+a25E4h1ZInqn8WTw7YPVNPkInNxmm0BLBBCBRvuuU
dwjek5bpuhygIYcTHZUFf8Q5Zmet+BxqTG5QWiPqOG+n8w4TYKQmYg5UjSyWaCBK7qkdp96ntY4A
ljabVTOupwI7tI3MP451by1WsRadH60hpG+fR44WxV2XpdpEhs5HF3hizR1m+QWkXthd+Vwp1KMA
dDMo5VzKMGVADsQteNgPIUe+VR1W/10qF4Ego6pkjiFg64JZtpSpki9DH6NB6RGzyWprkjeFcFMm
B98l/5OuYU2UEq7uydb8EgiroxeDZsC5AB57wcJstFXRMIAow/jHF5redasD1KpSIkwcTdUi+dqR
VUC/NB2aqLhhxiDxnNVR7kmGB989QRfrtgWFG8pxC1vd97QgC/l+ykJH1IhU35GCQYX4NVcm4mKe
xs1so2qLDZXAbFD/qRpr/CGKtK48/DVU/1cKClj6wSPSUoh+GPoDA/v/Xhcr7G4x0+eMVtboioh3
44jFGEq4u0v9yix//w1y2G6TQ2taQBGFDoUu45W7s7JA67j+M51V/FNtXsRXF8h/dCGvjScltmhc
YJHy45UN2tjftkhXnyz8HLha6hPzbyxkUGEfxHsaQhCGDPb5WmH0Ey+sR7dsSPvK11BOSvQgMTEk
lVrJHp/138LiQTi4C2CYpUKg11W368BRgJsRvKQkyjg8DJ2ecIvDWdc5ulCeIw+ti/dkzHOGuESe
5GJrIr7rKH3dBCn3TUvk9nfIG9spranhH/XzVWJI8leHRYX61K+ah3Ry/xTfU2sSQ6TSjRxm6mmY
RiISDN7P94LBF4OdQF05o6L8QrJVM2z9vQeWzQ8yjAZiYuW9RgrI2XAYjhZ3V7TphJD78lFSU7dk
TyD1ITf8cbHVuHKe1kkrll8zI9JkM0ueRzCtAa5suXr4t1o27j949gdsKNxuB1Fai8xSmeu3c8ee
QXWqP5iSqXBbDEIqxob9/R1YKjoP4im6+Y5KKIoIEluwb7zisgEhMqQlLh95uyCAcfaiQzyORPdv
dT/gmQgtMtgQ6rgvYsndObij/GCkfJ4CccNccoYBCCc4TjUHiNLuVBzOaoyKKNLrpwhkuUERKSQQ
/fCon24NjivCcGL3eRlfQYy+96/KouBrYaFacs0UQ9RoiZMzoFg0+7KVcOfB8UZrLLiHjV9U6Q83
s6fTbGVXTaTZ/vC06eU8tnXazt8ijyELZlls7LY29/rGbskZtWVkuXzEzde2kQ3ufToBykINnBRR
YFaneLAmt3JEX9cdL6oU86ZdK2OPi5lA4tPr1R/lTYC75eSteuU52Tf6RH8KOFc8r8kBw9W+y3em
MeMVHPotHULi5NfKs7uqaNIUbsvhYpSE4km4kDtR82CF6+u1iJeADEHLDTNdctva/vdjHBjqjD2H
yZ1OoLD80UfT+Zt6ECFfkPK+zPlZJMRmjc4V0/USeeJxg8jkD8zjrSTMltPHJ2VYuHzgF5TgtmPF
zvq12qZl2k3p0+BOZnSirAQXYWFk0yCuZlcR6l6+B5URmBB7rBH+TXWebMv1PoS0lRrDtNf2Dtgf
8DMCT2Cnmn4Ta5KRIR+EY7dn8OhBsbB9suupOlKvoZDuFbFhFDd0afsSwOKe1yUeye/LWwY6Y1Is
W0FoASsSaKygU8/4Yh0BcZoufgtJCitTOyvUmldYfpuRuC4W4hPOiDsrJih3qNH5dVCSQtI+H1zE
rJiiV14SX6rcpBW5RzC9/FPg4qzRFXenq25xz8MU29+wn0xp5ETRHVT5KfM3LBHlWHNhkKRl0Q9+
HX8cKi+6OzrdIBnLg53iT0jW6uvmhFnpZUz9k7KFQZuQo39tjO+W6yZkk7XWNI226wUJkHlUvcp/
YxEVFtpZPvrzttq0B1jkUXpl6okdKHqnsHGCnDiqdyzobxdxZAT5ZoLqpldB9pPXmxFi3DMhXyQC
LEZ8uUBE0mhXvx6EYu39AF1EDXU1f/qn0Ej/ANIpE8DEP78q5P49sMW+oJKPm/cWNSajKxS2ePCi
zXt9oX+eTqp7RHEkVmR8PU3FxFxp4Bm3FQ/qpSlOXgwFeSgxyx3MX3erRF/lO1W5Dx9qSP2oL+yh
k57exLtlcDPSmEBcfh+8W+Z4vtWWjNAaOKHCHB88PcrTMsvJUzAKcX8+FhoPMap3fcEvNZp7dLHE
4Sicc7GYIh8Qc3Qk6Uy3HMM8ypMWYLtlEldg51TMj1IBWmLOOF8pBwptwLrD96cOR/p5JYuhevtY
7ogdN4RUS1rs73NmNaXCDzx1ymxWhh6RzLBTF4sSMnsPpmK8I5PgrWBz6kEx14PP1PG6JuG1lYN2
P88ElWfBIW9UT8/tFqBU1k1/lK+y7QyX5SQfo3ulZpmlEfXLcipADh5OiRyZcN8OXf0bblqKuE4/
FqoDJuXd6d/QYzLE1WXnGAl7qglQ1B0a6rpUETPLzdepU78MmT4s30GWjiB3EgRE89GEh4eG3iwO
B/reryVorNS2aWK3p1N6tYLB+7P8Cld+ldx7bGyVnCV5kB8lwKGpxZOJ9jRXt+dekAct3gwtLEoh
bACTf4WiKZl9J5ESDfL6jWxVfANQjiSFAOMkRXVHKUwHtT1Ax21iHtfeGR2r7kCpFdwRea4NYiFn
2xIIfXAV/2J6CzHOMY4r9i2Yj4aWhcRLnwTzqn2h0Ueh25i/kGw4xhiPOqGsubEuB+kAkHK+OZMq
b3HShvFTqYY7cubjrneaTzQDcWZUmANbPGpaK5YvKSkAV+XfSTdLmzBeWT84T+mYO4x7blCgj17B
ALzz/GsLWo+9kgdjYLBGVJKREbkaWaLLeCEtFvw3mLBYBMBEkNQx1CsmQsZN3uFWXD8z5G/2gt1k
hKOmI+g7DGG3y0jEzuJOg/5JPiuxL9DNLeEFXJvNh0BMUum7tsvI/uwxcrsLEBFbfoULWzELyBw7
fHC8NgOBxhYx3lS4MP2bH8PhegGboR8MKxrDiOhNtyz3BO2O55DnjpnRWftobjdr5AOqYUU++UQY
yKwnf7jnsRmyMJliglue8MEvzGd5DUhQpwOY8IMEGXq2pyD9AS7JEn9zE6AXZ8Er4Qfys0AazXus
iBcEvOjdgf2lIShNkuycj6yeVgOavcKNRlnbgxrnHuQBWtIggW7iGzyrF56G7wgposO3WzDzIJTx
B681WozEKT8qI836xYOODZ8NqIR9+XZ0s+8vs/JppWF8lWnE0jr2emPGZYEejf0R4/SoDWJ+2VOs
REQV/maWoOekzAETvdAPMspNijxYwt7sXp7VeDvaW2Hl1JYr+Ln0y+xtOeHE3nFa3I9U+S8Q/QRZ
s6veTBv6yfahXsMhheCF3zlAq9mvRfwG4woYpr8++9A6Q2jFDVNEojXMiECPGsfutLoPidu0T2LW
1UyVpDiAe1m5NIsVpiJtp6PaWbjJ77cWpDFQ6YBuBQzXtA8ZTPyH1fnW+gkz3hbHk13i0TQXrGtg
4V4B3jFQrGvJ7WSrzdjqAmdZusREAZNeTB//gw8ZRXi/aQiaiLsTN79IY4S5fANsLINpkXWXKSBH
KcWjQdTcBl1FZ1DZrWY4xCeWVqvk6yeomLts7qIQtz+Qo7BmSJzwTF4wj3UeWFbjq1J5gii7DgLB
5V+kKEAD/TxDECXsB1bWqHKApvT22RKRCxS0V2DFyWUylXcGW2vwYj7K6SFk3p9DWqfWJKJ6j3Oa
FupEBRBt/poY008COQBx7lRVc/DtJzL8hUruI/fQ0c+WjXHfh5HTGrZPhktHAprYgcDqOML7Anc+
G2pcNUUcV8zNM7twDsC4oH/p/VQQWFuklqjLEABO8TxWhegHF4EgW0bVhAm9C8BZafotcTR7NE+K
H4UrRthX6TqpqL4AZM9HsDb1rfQDI/FLPlZV9Xieu87Bavl5WoRbmTZyldESl4QJL6op4ks4rh5Q
hEV6jbeYsZ1kSg5sdK/I/gDmdRO2tgAHfH4lOdLKX7XOPNoaK8NKQvlTo8vHUCwm4drypNg6tG24
x0AyJz++FHXE9vZf9O53n/fxPm2XQTLn5VqEO6XMPQSgNWalV+YS58MfiVPhdL09b9VMJtYXGy5a
AxfUjrQxVgxO9gTd9eW5xC82MeCYO8rF2CeRYkUnW80mVpSAKamUAziHrRZkEMiqbU0bev9Ea0kd
pgeYiEZpWcczcg/rUXwKELC++PLjxl0fT/v4NPlO29m9TUXSaulRLbFmejcR4i2IaTljDZP5nmY9
f6yckETL1bodP02GeZ5wQa3t1U0XEniCmeRTZm2qzD9KgJspRfDal0MjA2qGlolKxG9+3MuFHArg
2D1oo9F8ofeQ+qTqhfcx7Vem2hk8B4VlKW11j2Zc9yvEIC1aQhW/goHbs2C3KSziCEm/7xE9yscx
Lg3t/ZLZ0MUesG5IAL2xFBTOpctXuvYBBAef8DHX58IoZr1LMlnKVPMSfo7OgfW+ft4b08z+kVRP
Izk77tuAr+AqgCJbM71Wbl6g887flvjfKBUji1BJVKUfLwReTcBXOmjd5UOUiIAPut8UQRgHQfQr
2K8P4deNKWKbuFH+qGhDrLyo0Ex2qiciJ5Bvi5xFghjOXL/NTETuAPEz9tJbCBQTldPw11tM8Z38
yEIYHLodhL7OU2aWhFo+JV34KHmsKPLBt3aZgg8P1lb+y1aqOhAOKufoIJXrOCs7bRDd14hUrB/b
Y14qk6BX1yjF117o+/rgrE72HoGnscy8meF0Cu2wvnEL3gO1BwQFjdmeJUS8+f06TRmspN5/J154
aQMgS8Y0S46EhXwe7L38BQyz3/JNgnZYzzwojkg7fxwQYKGLCSmqdZgVdGNp/bzQW5jLjzOgy+oz
cHb12Se075A94gHz/SBOoAo7M3z5iyErbKKifULNxH4vQFsA4chcrRfWwlKRggjQXppIZnIf9GiI
WdgNj2Nmjh9HyhrLinxeIU9U3GS+I8icIlQwNRllaGeuW8lHf/qn+GrirftaHwJgIh1V4ff9i50A
vUQzrkb4GeAauVP74mrsW5FUdIPJWGHx7mHPTehaOYXIFcpitE24o95QWCNn94/i2HjG9nPj58cU
7xUnE0vVz/IpM8Gto4h/62aYRoXj/84Zy4O31aGdbYKh4Ap/DaL6CgAHiL4tS3h6M83b+8H3fWQ0
RYTlgm2J3kzHZPgT76iWC3MeFCWSc3b+EnZ2lSPAHZ6XmOVwlPLOcWJtFGe9P0RLXDYKFXXWF3Lx
rHD4wiCicGy3yE7c+fbq2pxFDlAwmUH5KOPO1GoTFhsvOs++4xnyOdP/HGBGgkAgbewrljAEkcO9
TBJjLsVKabu6ZXz+BB+lueACAHdtr/e3DRaLchMDmb6qYTCqMSlHuuz2GKna0ulf/efMePLElK0N
oQ/CV9satML8uW53ZgXdRE9DvUKeVEnZQgBZoBDAUnIqfFhVuEWkBkwQpuBbCvaqx8IHNb4atO+7
29nGhs6TKbc+CqSzKbkLUTMqy91zT2Ulph1iPS8bIhAVYkJG2Jz6ATW8x5R/p4cEs1rPRFf8CSrZ
YKmK4o27laxBJhu96hyzf9XFsi7T/TMPx+xq3yWXig6egCI+rWJI7Wtztlj/vMDmBVbayzy677UL
RH4/vYc43YlnI4CRjn3LkBDlSkTHkZIp4w4f0v/9FQVMjVzF8UKtcLerNKvzMcg4D/snUL2ARfbz
9A/nayoeeQlwi0CHapmNaB+517wMe6oJ4U9CTmcLWOubHO9M54WcIWixP1ZzcddEhFJuoung6MDt
0PGjNt+BSMNvQVrKlWbT2vxgPZSAgNbyXcHKHvQR6NyssIe3vWXqM6Lf69SXeZffotAslqRBYE6I
rOAPO6q3FB1GGSlP5bd4z+LTEmDcVAwT0yHOXHRo5yvnthjwdDIXChbnEUZSWiKqJtV162DLHXkf
aGGHffjybF4mKxpvjHpMc7tzBD6cDUBFPVgcUjggv07clGfVFxxqKnt00z0zBjpVfZ3Sanyhp/Te
K88n7p8NkmYPBOk8AEhGLwN5ZsCIPlabRYpVsxcyAqwovCC5O2+5RgeXt4fbTv0rdgZoPf5h8fuY
wzXM+Pm3A7aZYix8E7twb3XNM0WYZzlsDcOK1ACYB9FsI/Mx0my1l1mI4qrkgmpP7mcOzO+qNnQ6
9ts0RinPElQW5uUlH7HdjB0L2S2Kju+KkjuiNUiOxd5awTbrwg2ZTocsOuwvHHjckkLY2p5RZhUs
9eKvBH1vyycjHuVPRSauMUE2rP/Oec8VnebZ7vc309My0qJ40bkLxC4DP3FjyeMD1b/9gLiH8/sg
tXI9pFOrr45mLpk+owoKkKfkrqusTuziRWROy5Bk6/T8Ij8NhT2YQ9PcgWnUp0U5inzo66JMbUuB
gKaDLcDpKeJChlUflw4uJOpHfe0Q3DkXzW9r4B8+WVVaK/q+c6QVuQU4lgzvAOnaS3iSU1ddMaiO
fxTMxNpyS3kNN1NwZ6ZwwGu6Ikr7yGQzjwtDLMaoSkxwnWzmYJqyigllC3EP3qvmOjJ+Taagyha1
hV4vzTUZAkwZYi80AbQFx9y0dhjmX+z11C8ABeGeh99m2TerjPoaPT3sSflWDPF1QAIsLb8gz31X
Zn2CSHA2axGpo3AvZ8+COvlbgbkWBvGw1q/UpnyGtXwkrWREAbu1/znr1dVBn3GjbymjImwlBt0g
VvMaRxhhCebzgO4QAbdIQTfcRZwJQL5+5uB95yhIaJAafKZyd1lrNKTAzgH4nfDsGtrYt5u50ezk
QTBbAjXq8rrTEFg2r64TBto9pXjUWvb7gtTEAABmesh+J1TpzeLEu7ZQIBXIVl0qSYK5jSggutrZ
26Hyn+/MmSzLWW5SnHt+uN0w/ZfhEUVXjaS4shF+bSuOgJ4314gY95m6BFGO51OCkrRlCH19ndLX
LJvXYdwm9fwm6xYrCWR3HHUPmRhYEoPeLpcz+e7UpqaWYJI5zEyYySTtB52+GVLZlksdVFhGpfWh
jiOVqfvyjtdhsBhVX30Mf9zkcM0l/nFqW9oIegVcV6zKB6rIfC3GOomm2qSQRoXsnPuXc6A+W+Qo
lGYVvbsQdFFWGuQdsgfNFJTYPtumH8BuN/yWwHBorxA4r6Xa2pFNOUgBDnSfUhKues9+OAZFbUq9
hyYXJmi54uYI0psyUUxzP51sXPxWAxuCuWzCOfsA/9zbufWsbwS+s73GxDasD7AlpPvgzmxoBzpn
dzOjlhXTyMI+3cWTk9y0olPYRD7JEjm9BEFcLobk0yY+WqN1zBo1V0jaYnNfQ2f8ZKadz3HttZhV
sSVEjzTftQpfj8/hF/5VsbFH3MHaSwtsu/CwQF8tbvSwTgH57L3XXaj+7P/eq5AVOKAc2ZyEb0zi
PJrI8yn6p90qDA8urgSD4S6zThHaSjVaGuSfFErQntjHHQOqG5IkV45EiF1DDNPInZy7yCn+Hw0G
hA0JZt+7G+pgz0QoZGymTfQROkiIwN34KOXHpwFLGPzThlOeR/B7F6VEl+vRkEzUYlW4Cc+3JMYR
bV2bqEh9443uAzk0l3VHTdOw+mIs7DHQiT5iuZyXibeDBl6CK2yiWKxvmz8msg+f4MJI0vB5s2AK
B3vQfrSKtjUr3MX5uinx1vygFoyojFkVOd1GeASAbCtMTNw4h1kgi5v0vjRW3NiUW2G2yFF1ArEU
Zu/iyQRpRHwTcbw/L9P6cfQ5ZSmJFPtPD1UfG1uzKk8tCj4Vs5B8NGSqftqbKmjfegEaIC/wwNXu
mVQ6NHGjxE0xJl2bIlQNOxw0x879DGnQXZs5dyhD/oq6Kp6KtIAc0cFQwnAhifr3XtZGcOCWBzdv
uMHwVkS6Iwl8qmw+7TdA/i6DEKZwND0f0rk2g6d8EqHZcuVyn7vC5rLwDPKKDRz1MheDL6S/4Dil
Hu9pQ2ubooZOSbHSpj0aUxKumtep7Kpt649dT2RMKKpRjzTPfR5NhX4eh7lUMY+Vt4naLUEIl4v7
jHeLqN8LxX5ES0x0g2sbjaUKjTzfh6WdQMwZz5qDez6ZzeV/WGmf9k/vOZ4wviv3PQCvH5Y33bNs
u3aFOKuQoUeygbHYAH60mzt7p2YwBJRi1bh5kde8jVoU4ZvfEVWirhpMCHVWknHcMhEscxkGYuyz
NiE35vWlrScZmMcLJ4MrrxtpR9N54iSbKR2+bNOkTr6y3gHprZGD/3nU/EMMnHXbK3QfqZ3pGgiL
QQ2YkZqXA2AT17cgEeUWqYe6IBRTynBVKpkru2ySazqENyAMGZ1QxuMSIS3fZ1mvNP48vmGID1Ua
/81KOGBXuF+MX/kcOKTrvsFrL21OIi721BC0eq4ce6mHGKjTSG7j9khWdM8lRJXD6qL0TSn2RbUz
gWP00syAcV4h2Ldh2LP7e4ExyN7tI6tpzNMA3fTcLhYcya6yVUI5Jo+YbjD6N8hzqgM2U/03U/QW
/Ykn3C6lRlYHR3+LKWQQfzNFEsVYv6t4FEPoidsX7b4EoVA4jgrY4AC0t41NnRanU56dt7671ekm
pWhyxqStF2FtODoaL9DxSlxuNOcx+aNxY6kl5tF6uv5v/ipoCjSy52RhrAdm9NhGAM1Y1d5ME6iH
TP5KwhMRMoWTmddkXFyWXZFXlEp7dmi3K8gKSq9T5zBuF8jEDgO/sUq2eXHa9nVQG8E/iaT0+WoZ
F85nxZTaeJeuRMVJCBfV0I5ANtn0ky7QtmwVrZirpHS9oL3tmSuhdLsPCjOKC7Bzr7Qy6sqc9uzd
ehBZKM9PzKPQ/c9gIiDPvB8Jll+jKjad151/e2zxehNKiF8yjVRT/Thh+cYltVjWCgqwj/4OrtbX
VHCBiMfqOdF2jbQvyKWESpPofkjjAX3Ax7VfzaND0L0QzqAZ9/KdD5TBFf1ytHDUJu6Yp3j0xS8T
ruiyCodIgTGxrTtImiaiWP2qOuzpzkyGTemvbV3tCyghgxKUYUjbhCyS9GK+bSSXBnRSlatFhKo6
uex2zkosM3YjHwl/2jIB31SX0I4cq+ADKhBVYgg1aB406gkFAQDi85h+IcMrxKPLXaYjh7WofNhn
GdyHew5Q/S73jxtpbun55GtB4DIClrXIbqjNJwrO7SKiOFKX4phAeu8/rP4iJcH0FQoktPY4VB+E
EFTC2TqSR2iSDjZbVUHw6Z9ef90wqeNHWkolhhOqcVCF0uwJpvdHvkdYhK3geKM899dZJNVLoL/a
K17dnh5P5HMWxVkKw+UO6Yx9lQLuYo0OOdtBa8SiO2MMNfDxl9Ym5Fqp0jWuKeKXkpyRBSDmRMz9
4ztVfqbPoubX5lgRHMDn9p2Ws6ICY9ErdxCRd9Pq0fs7LfLw2MeMbeHsVMwOcJTgUePJwFkDG/2w
sY7XjHLvp93ococPjBGB6WohTPIoRn6sfcwwq6p7Q8HxUNmer4p5uKvYjI3T/6izmpJ2X7JqTS/K
84/0lt1s/mkv09LgqgQGyqsQdmKoLEsgl77M5FBJj1UOMCZ0tFdNp8tJBM0vZ6Q3v4sBT30UQRok
DFmAyiSBT98iB8I1JAyoxR7JQnDaghWG1VRLYROWNGabOv07x0UgWJHDRvIVrs4oU+s+aSPVEzmW
i2HP9Iqjq+UFC77vNSpEaJ/aQrr0lNFtyeopT4Fn5UzOu7i8zuEXvMdYXsm2gysHFVgcV5YGJvRa
yv1hFb0v9ElwtswbJCMwP5aG55O6QQ3iEvqMGlhCKFG2V4tabDDEYqWupOlVoWtNpmMyiMinJY1t
8i3rw2OlYJPSza/HypMsPrDzBQpyvZHvDydnQxEf9lXtfyKXZGXJQMkE74a2l3KRkQ9Pjladb6S+
NoTPCZZo8WX0ame1RzQKSuWSV5PXZbhT9HL3sE5PvYWqfND2ME7cuQLg42vBuD36cO/voYeMbtuw
zgpl/GrNK3BciPYPrRPMyxYDqHhrH4KRh7jJM0q85q/lLNOwezbpHg+a/WPlj/5qM9zZGNbB4qtd
klHvRH7cxOOU5JJ7KE+0/ZqnNZsTRw7BwxWEz4R4dweiarXuSlCvvtL4dk0OdA3iVt8Eg9HRNHt8
YcaE+qQqdQwePeZ6ax9ab/nY21Mzjn/+RW3Ku+doq2eLu6SX0R6+UK9Kk2bxMXJm9gogFJWeBmZ7
YS7SMJPcxeeOROxMKb7dzw171u7iAU9oHwgFmCiEx9fbkWowmuHEBVNKqziSjiuJBJG9AjI/TJbC
h+6HQ6Ect1+gVq/WWW4vZal1tmY1tRhSaGnCbv3kLLBx1VzmxVx/u4M4ezhH2lGfCfNENGcYmqkZ
hzTMnG9Ov2TX5GSbZdhHZ0NsB7JSZjNhZJRP64RZkLjlGEI+lG9ZkV18AQ9lwinXfNPHi/f1lYtT
zml/RXxrMLCHMUEI2Ba3AIOJP+aPoZwuLiYozbzMZByAjIKPbOZuYhlFZ66Bjl6QUZkJAKIjNNW7
iMpix1UbAcmIacHTHCUZbiSXeQLt04mbeht2WovkECwMaaBHfjetk0KN4OUz3AoAT6n6v7/xHCTY
GU2CjvL9vE554tNZavbN3Hd/t+4pDfb7/QeQE033bbWKslcu5Hq2puDGYJjSKveStp3+OQMAU/K6
7+xbJOHjVzM9lo8F8DDwt+QHcqN/NwNZX/B2VE9c3O56FwIXq0AEz6YQwF3N7IHTwO8I49IiEA9K
fWmlvSfOcLHJx05pgimyAt2N7YKH6pwFVWo6KysRJ9YipDeeaEHwYpfOxu6B33GKEBURDWS6+gDC
w4wM+aiWT2VXXc06XZy238VwiY8XjVevzNfiTG+1EGYsX3IiRCB84xDEvuOvadQYBFFuT62wtg77
AYoUdnRRvSnckhts714uLJ+jb5kyvHIMSh8KqS6Zo28XbrNvtd70Y/IsIgUKIchQ5Xs0XWn34Lyb
tZDMEw0PvU0clfOYiD2YRq+BVgXrroZeW6si5CmI9mAT72o1RxTFfKtsnO2q8V3S/Jj9iJLzMDwP
G3YpXQu5tugtRAYFbf+zhJYp6pjjNuVGKTSXipBf03O+WxoodyKJW3qI4Bf0mfatGLS0PFibANhA
km6ZcNwHyyhFIk/JbUyma0IKeONB+M+bDvvUXq6eoJJEXEOn/GIGYBstELfZ9GohidjocyU4w4rE
msyTvscRAPtAF4xRjuNGs6dY7dyjS07WdcpnmPvHpgPafBTaHLbKNvrbY1fHL0XiL3cHqODXsn2H
wAZux4x80u2zt0KMqbUqKwSYeHkR2Oa+ED7Hxx/wTFyxZky4F79D6Dqo0ReyZE5ZGeZPfyWrVP9b
bvXzV0uTk32/546VbZbMGFGl+NVFzooyDmAv3TQ0rLQrw4s/5+LAeQPTTFMyzNmoFBM3VlavlsRp
5RSbVBbFoBWKEghb4WsvrdDfpaA1ZqBXpcsaMj/yzGQymxVY+CJJexyI5+edJc1qmTmJ9cENsvFJ
suPu7mzD4P3/olzujUcidtfEy0yccrTcgsgIsXP29FXzIyqvbbhQFg0HrQERkMMQZh9Fg10uhwp4
ZM13rgjof/K1+Q0IDXHSvDLSCGRcCTFT0W89ZiQYmRw1V9uIf3yMnbWoXWAva0YH7tJ+touChoBM
QcXw1Je0vt/Lc+ZZSUqHCW1LrH4ktM6TRrLNQy0bdu55EonYkvtbyAkBsex19oxzDAj1Rhhi7Kk6
qyPgej3MLPNXTqHxdvHIwAXDAAQM4mxMNBLmcNTl77Pda+dM/mj318QjJOCQ/IOX9EwOEgAKQOWn
hh0/9H7bB9PFfhhH8wU9knMIWFJOf4bQJSkAMu9JxtshbJ7wzywRZUbX9VD4CEL577VNnf5kDS2s
KQKF8/+yB91nMniOAnYhfQ34A7NMdmUsX+bt14AGC0GGt2fFPNie6AGDoNaMrSAwadOz7C+WaqE+
FOz/72+EDh+e+2crhmdyvz8Wvq6RzfMl5wgoUI7Wucl1gdZBPN045jM5fZSAZv0v0PeYQFCW5a7u
fOd6lJwF/liFD9HcoI3Schl8e2xBVHdmrJs0qEWjDZPiukdIJjfbexGvHMPnbDq0Fjd82HH+q1sZ
rhEdOzaHD7DojT8XwWs0SBg/lBoHVw7Bu0aTSQaQoidajidRcFJLZwyfWiNu/QXCbyK/1XyRBUMq
XtKkww306Dpw65iZZevfPPBpjABq3Rr4cYEMxjMOpU6KFp7eUiE4BstMnDnFyGas6ElbAq0gX3Ha
br5C64eFQZiTPeIrieldZPWGycRiRt3tvazlgkIr06MNXOjVZaAJKT3Wnl0isSdby6ICvMmh8qHx
h2moGbvsMm7xtW+crDms1faeNAMxmwxIcK3Y+0p7wYnHPsK96KBwTki0ymo9WNhlqZJvvcL3YtRx
VrweKGAKdGFFYh15Bcoegmh2k3VY25ipxDjw3iwVkl3+xERfDNxgOpU/DOWX9VB9y6rBdIgR6miB
SpCrilvI0YjCEYaW4zQaQ9/kpdKFvUGRi/2lv2GFuqMx3f5abd9m/+voyj1BKuA5+5IhOCwg6bUu
y3qS4rpKYwvykXDl1HvR8UacsKYkKvM0mVqyKHIIsHCJObwB+fPDgh60ciuZDrz0ihBel3Q+Yyt/
QNPILqVOcgrt3kkPhM1pggYvhZWtUwiNMXSA2A13TV+XsVO0oeAQSvpJz9M2hWrw3FGjPcp+u6yP
Jhmz4aUzAvLb/106z6WzBbN42wKh+cjfFJdDeu6lx9qKO3gZzGuiUOIsePDNH5QFnKhO+B53gwSD
Z/4UwnOXrpOWTW7NmvGHQOZ8KoQyt7LHWXwcrxa3QcfNsvJiMZKNo8/Iranov3huN5SPz2GeAuS7
+2h9DA4ard9BU+vXFAWYMjyZNALSZ/u1fgbZZtgTaWI83Qv/hKWmHB5OiqtGWD8mf1fKKJMFjBZD
yHUWeCX/nD0xzfMJbphTycqs1fVJRoGnWkRFBs34PqyjBFGDpXbv8Y5jx92poT2JwxaVldk7Rmfz
uJNSLMXlvemquB8CYKLT9OfJV/QzqL0V2F+G0CIyo2f2WAxKCH7lzb06oNFywuCf4w6bXfQYG1Vr
4zgPWsWaeWejsEGwcNbAsHScCHO5ADCB/RQrzGSg+PGks0tvZFatmtC2z6Up2zmiQis7PIZihXNB
jN7Mc8daoz6S7ZZTTPM8pwHFVUzi1KFDDHX4JC47cJutBx9UuR196myqPfwAb27CtK9lda0bBVyZ
WAWiG6OAL+GRRBoBQvUS4EORZDjYdvqKxLxs2D9NS7Iii5/x+OLp1LOlfkbhhEgQmik5Xdu5rMTK
xNKwhSp3ZsK8OunM0QMSJ8PXGkjFSAhf8MA4uPavkK1GsuSiYhvD1yyd6PWH3malEQvMLH2U7/mI
rLUGfnXYAItkrBT4LVdLeCj89H7ydG+4a9a4ezXB9HhF7QTgY4+v+W4J05Y1xZ4TIARTbtDkqpFD
97VjY9adhKz0nG8SjMXQvwJF/Y1ZhdkKR1QhEzYJmpcgqLe8U+l9s/kVxKa2XaQdOGDOSvW2ds8J
IQm2YPzLJBRBG5INRp+VmNskoeUChGpZ8ox+zZiXg6Xx759KDsJfbYN+9qH5nRxWERcUwvLh11U7
aw2x/tSV7IEPq13d2WwgnasJp7OarGMSspDh8N/3Cnj9/XcZ0EHJqU/QvuEo4ynWk6qEETWCAEY+
yP6vr6XbEDAJ8ZpLoaOWlstBfY8e4L3gUJGsQ6A7BuBJWvXpERrlwqqNm7s5wINnvSxfRDrVm3MW
hgQ0LcQoQ+YNzrLTXA9DNuDxM4YbIVn4E24jLX4iOXAQweqLTt58b5SYfM6Kp9rr63vNS8M6OwrT
1+n5Q00YzSwsXfCBPgNbeeAvx+7StHwtGo9kGM41aM9udV0i4ckl7i0kws2Cck4h2kJpPXOk2DRn
wVd4rieZZXMymIaiO7cRldJs5eSBd5ZKo1Rx9SRMso8jVLJ8VATHrREPLIGr4Lq6qCKxJMPZTFrk
N47CbqnLiOAuA8RVo2IUm7txBU0gDndRyYcnipK4afKOx8VXHLuO5XiDv8GkqkXVJ5E11eSV/iA0
BtxB8wDCObW+vii19naX1qDMA9Jy5XYXsq7w9ns/UiNWp1+G9Zgqz+rnRqoBoeqlPsuJpS1uh5Gx
ZpAbOk2uZy6SiOK7KdgtiwIvYIVivZnXYbHCYi7K3Xw8JK/HoSTxWEUpkzb9q5MW1vaGl9CWpLmD
04prIimIvop9nwWiDpiZ+UpCql8zyXrK3saM6i5jXYHIfoISnb2xJfThr98lFc1hVvTwYGNnsZ4R
pPSn3LnrqoejmwOqk83miLCQrEo5yyGXa4488O39FBUchY6CDRuhVaVaGVA7gCeON5VjxruU1mdH
qRHAOfMv4s/G8n/TEoucBkqysDUNjrFYLv2yWon4PAR98hWm67ELf6cAJXhimP+vB0PkCq1zf2Bs
Id97LHDhhU64go0UGkkGP5EghmjimB6cb//4bzMvHVLTXyFAT32S7vYqql+pnr++pDf/976G66bx
t8ByPfvdHQnJROPWouta7T5FECKjzZXdLC6q936gs0TQAF8MsM2panCtYoynYkeGuBflgdZ0zyhl
4ImmRJ2PGZyMBq+IOg/LGJeGdDo0iV31s6LP3F4/SoMwGJzI7gvSk8NnSFQXqSVqw9OBItxmAGSC
6BuXVnb9v4wwAI5RF2X4+D/VmQzxERwZb2bRfU5ACve6y/tUBeN3vMKQTe3fxJkoFqiMXix4QZS1
bAuxSiiSHnllMfetjDpx6vBke7RKY3J4vPeSZAETOGEAOLUl6xeS2RpWDRS8bpUbKYhv3zNbLwYW
c54tMJpiVdaCRIBMk82eLzdw1kAx93mGr9UOWjiSAutPqpqA+rqd0dHe9SdnEbvGGhcxVM7ioen1
pZ0Z2VSzbxrtRX991guJLQMQFGJrDzjaohrqhscNJkOQytZ/ZOiZhMsZO3ozhIRZh6hoB1xLvuS1
sd2sNPc8x8pXhSFdqdT4oqIyHXHNvObPL3jpeDNlv14pqhGNujjQNm4SNCA7puI+IYXjHmv+VpTE
igEdYrxmIYvsDEX+jO00Jl/WRriFnHd52pjT9++LYWSLPuW/bE/mLjuD8Nv+IUzz1zm9opNi99H6
EpD0/yHkS8c1qOOrzUqRLg507+A9IW0Y8QTY5vklJlhULA9We7/Fan3puGnfhH5U5XrjcU7iUU50
SOlC4kGJ6T/sqE8Wt1zylcplRd0TmxV3lDfWeLAy4t6LvmkT4v0YQCalq5hdbNRB2QvwEsP9otWn
HvDESweZ3SMhvtBoU2KPEm880xWYcQwz2mkw8vbId0cJRnb7CYiRq4PSrxSLOEawQnYjugKIh72M
STIeuIVIj9UtZ5i25bSjX4/eJf9lBEmOH7nyLiZu1kiQC4TzSwlZ8+Ei6qMPKQvcYtsetXAV7l2o
uAZZeOYNu5mgAvgSfmTlE9YnS2DT1EhVcrQUbhDMsa1wwUbCseX9oLfiAvl7y/VkxBN+ZVHTSRM7
yJnzjCtYNeJs9vUKD29CQ/CP2KR3ayQSI9kXl+JrWDekWGa+kcXRZTMKmw5o2gWpNeIiOx3ZQG2n
bTpD9uozgWpSWHg8Rp3mepmToFSQ8KZ5F5BnXtQ2RgRNNeyIueYG3k/qbrD4xHXmFsF+8YY5KnQQ
z2yQbleX/Mla9KFv1SKIFpg4z69rGie/AAUClzoKyG4VY/irCveKncLnXRr0zSrJEPqG/DQGUYmO
a82zmdvQLQiJ0UBO8lknEZJQn0lGz+uIPkbOKDi9tuZ8YZkNzsx/ykTwlHS6pZJeDi1tfazhQTjH
er2LvhKDhYCKE9uMa4TUDRD8d1xncPczK4+21rj3kOtRRh/HBPfoGqeiT0YRO8lvT8BGx6+DpbdN
WhDchDNGthT9ABbAacIx1r2ZoWiWk7nC8FbD/ny6FGzL4c58p34cj72u8VJSySeAz638Rik68pUV
3fErf99rGprxCXo/iyywujoK1BxstjeeJcJlHOVa8I88+EGCvjvLCyAWV4fL/taTaDBOQ2lNQ2UA
a3xHuRwgCwGYdBrs8lOKeIIAG2vHkSgWDGoXde54O/cPhu8mnmhcLg1bdOc6EBnj7XRQqaJWC2EH
fND/WBnGPIwKFOfo6g/IMuwzE/zvjLxTevj5sdvv8L5/ymmdsUifbye8Z08dAdI8poV2oA7Rv3Nh
sonJbPl19ZBUWBZ1jEsL/eetSYIz+ZTyK46pOP1BFvRfOrxm3/y/bHk3iuweSQLtCCjDVZtYEBon
r2c4/Or/WApSObbIuWuCkkATy9robthK/tGRz9akrVXPa09CtUFn+e5cqMSVmkpyVBmhHBeT34QO
PAWJbCfzi/sYNpChCX8zh3L4B4EtQQgeKkzCqv13mduIJTmD75BQTc9GR5e/PiJfUyPWT/Zcaz3I
2ScdhhcYThKb0/k14YoqMZdUM8gOrHjyZiubvMrEPa60PvBUSzvi+2roIEP9P7cVFQ8N4YArEu95
EVPQGPy84Nzkl3khDWosKq874SeCfyYHhRILbc6C5lhnSSmnQoEM8y0iN4PeiAH38SmMmNjg5S/X
8MjiEelzmOc4hSFXrdNKUi3pz7vx/K3QOm1yBLm7w3iND4GHQIBa1/tz0sfUIhX4NBZlvyeLD00D
7L2a/6s5TQ+mTFyA3N4w5Ff6TzB0oUIU+hsWgSU2RA2gs+cw0Uyb33wusVYnX1sJoVOiEAtlOLXE
FYCBp6HiOuw6+A4tXNOBaUvURJTOIxTWezMilJyNjUSH6cIqwzaZnXZC1i057sQEX/s9ITa8mon/
lzpCJXX4AU4U7Moymfdst9dN4CWFQVN1Dz2vUhZNPt45k2zXpZsCUw3XkUZ5hARtfNEu2KFkVjYk
CyghQfnYYDYVOqn8jMVFwdrFcJ6DkvofjyfgOFKMas6GIgz9QCNG7DIuiC8/k3HJS8nyUIaibBNW
nS1NkGZ2jP4PyhdwYkWJrJojtegKiZAlPJPsigYcV+NeNQNXaaNkC6tyQmWTudJOvts6+DCOOQ04
yCqW825l6QaYgpGNw7NAaIrUzsPoYBmNvvZL1WA+P4P4yqTMPpRSwLoo76VpjK2s7X/mYQAxtxg3
igi3ZvTXF6ULUziXaABVxOG3c7PIauPuk19WwATyggFVRvrkzQKK/AgFR6yMJjgcXkRPqfW75NJr
9PeeJy48RUHrlzTui4vFJOaZ4mx7fm/PdjtgbHQhWuVxkfiVM7QdG8Qe/EOLzSm6NIupBOjIJ7i2
D7h8dPED8JURRh5H371ik2/s/A5ldxdisdgv0sFYV2ffJULCH/ZzTY/oj+oPGROwzxtuNiJkm9wI
oWqMVxJ6H54OGh2qLTC1UQccqbeyK44uj1ZDDeX7ktsjuQ3jpROOmkR7LLOQQ0bYgwRb/M8HVm2A
hnrFKvQPERe20aM8ELilBwBdVKUOOKWBxAXBo6d7JZEKRoVnt3twJiWyMeb/X1Yn5rcceDeJMe69
pPV+mLYmA9WL9lGpBlpWyxFq8G21H3rabqpquYvasQPzYiGzLQF6ZqicOEgEAKrRU4+8dtmFN9JO
KOqtXd3Agv/NJe9B44cK4Z0wDcfFEEujWvx7rDSgnJMviYI3jkno4SnbrOXo1HaCwyRBgTZGPtnD
HOwRMlv4IYkH3iYrwDr5fYW7Bj2iZiY79y3bh7x4c9ZjKJ6UmZQxVFe6LzPqIXesXP/sQhNszJB8
EQ2ss5b1rtD1WQPJ72HgqHRf8HIsbgulE9uVT2bPOLQugBe6lWHwObrhDBPSLG+JCFiUiZLx/m+x
nGWk4s4iUzgandaUqoJ6AXE/dX1ZhZ3m17pbotNJyGDyTH0tUpI7VCJpIz0I07FFI4tflLDNcDji
KaISmyTeRp8i3wLfzYdLAhcF29YgBckPnYbENkLTb+PvyRNqobiRy4XWsb7Ml8e4cSoYTqA0SBin
Sw15Z/6BTkr3HkU0WzChcbOxAtifsJ+9U7yeWnOAmrry0iAAynuZNwRMVBO1NFd55mL08bEXnjnM
ZfbWrkw5kAllbpTdq2l8L/cvxF4AxqDX1ucqNOn/XMyDdMl6MK/71a8qUL13Tt2uEb7KWCPFMDE2
/az9SwPeeuY9CheTLnqTzlHLueCbHJbLwvFGBYefiRQh73Y316wdhYVV9czIqH08Yb+WPUXoT20G
WQeWxgMfTWa7HYTDqSAp5PvD6yTrkEMW/x6VXlpKVulxKqmmscQyBgHcBiWVsbr9FW1gFXafkK1C
GYETa5okEpkS0pJC+84PmhbpjnxD7a38GKF9L1rnsE6me7jHI1mlZRU9LGzSB1mZsh46NT3U7lLA
hooHXzG4iMOaiHXyaMs9d8f9wkPqptFMJ+CS2ryuMlAC0WJ41MiiVgAqMlEcGNYof1XJ7CxgjIJE
ShKdPSkYf6xXVbc6IXiv6d2BEvm09M0/SfTtgIaUFyRJg84JZYMjQSm03iltf834kb8RHQhoTf0J
VzgEuZAfOY2j1chbtjdtGJyrA6Ud1VcWwwje/mm7QGKIiCoPVdpETsGT3LXPxhIfLpARv4x/7b/n
7nnG2yonyWb5kvNYkUM6kS+13pXcPlZ42+EFAZwptW1xKXU3uVJ5wMBcTmR8rDsZQRctVON38/F+
nzDCd+ei61evKP7KCfmK1B/0VDsga9m7iFJt8N6MGy1vqokH7eWWEcYjRHuIhX0GxbgqSppXf5I/
rmryYmn+F4gmyVRWXiMQoPKDAbs2aCNGGEHZvUtNOxMA8LkZmG3EPgUJEd8w8KgbPZhqNaAKZuzP
o0ZwCsqKSDffSNAgJ34wR1KBRRNu4W3UUItSCEyNYVyB447nL4R3WfmcVZdn8ZQey+GM+anTL9r8
/WzPZduz4l3GlJ/E6JPteIi79x5C1/JHJYqubc+wCY+6mqn4XoqED0i2t+hlrbPaJC+DzHgph+0D
aULhxJGLtqlDVhAbSACKdUFbQutbGV1tllDLWfi07/g4rgCuLO2XB4RK+a/Yhji88PpWqKrisc58
9ucCD7NRyZo1z3VvhztLOkI16ycohekIQa52pdk4zrieSBRKQxlvXuKec++tI963pL45eJI4cDnv
1eDy9T30Eyc5MPqiflrWQiTudLB0Nhnz0ZkVb/L6Va8tYCquaQVOjKAeoZRl0Zanugn2yb6as2rF
85on5eGsmIRN9qdnk9AZ2ueEC6VXy9lFx0FGAqMOuwKhgMvammBLNghvKm7GHq461JDJGdz6DhJl
7bW4WiBvfgHTXodi9Xq5HpbPNZyfRPtYu+KIzcDkB1VUfWM4GeoLC7CgV7Rj8t/vVeKZyigEi0n8
XMGGn9Zar8JW9r2s2amIoc5sVBVZo59eBbKgYnAGUPhGRLjfOTzbozjiBB3uIondrI8+8lWm6EqC
qA+HGwWSTF++MioSCjm8nsbjLIn+sYLYw2jW4bXOu3RJRWarfOJwpwchwiMAOR+0LXebkZfLh/YD
ZAZZPRC+3SkQa+moC3OZR69aFRFNoFu37ilgrbhL0DYAJSsbrIOjSPN+LcLOnhJ3p4y4FQ0RaD7Z
iR+8cqXqhpCzL85DUznWrD+pVQ8UyfNIiMehAn/Kv69MImBOnlr+hMYENbSbg0I5Qxj3D8PPm6y3
LOSROQJAnKFe1ZxvJuUv+8KHkWRYeytZq8SSE5DRd2l4tS63B/e5CPmZVTMNcoukbCiyK4brxH5p
1NUChxFMhkB5tfgfCGgf77r3zrnxb6dJcBTajPxuzceTaAUVFD37SAsmP1qNqTFT8kq4oTeWdU7V
pwIIINjdvFiSAqr8Dc7S41y4egO06a5Cx+31h3TCBcGfBlgwP+1QimvmVqLMcUX+D7E6DgGGq40+
BL+UhyyYJ+asqSf+Ruxwo9Bnc7kJjg0dEUzWQcsoQPCkhk4q5DcHvCDICp22ppZcY6YGtorAW4MO
lw+LFkFwNCE5pbwH2B7L0LFdPRcPl4Lbw8/Ni0NGywlefA/ivsPKaAevEqkRBCBVi6U09Z83ZLdb
7MrdpqhjeArFuh/Chm1Im+rTLCb/cDN3WrCMcbreRgiHlQxGH+zgDJmu7ThT5qCeW+AA2Lp+7JwL
r37Z2Og6xU+oBqqMeS06Mmd9xmlEyq74IyqPbtZwOfLgcx7Uf3Cdpd9TZFrGXzXqYPcuNxYtb8uO
U1PDA88UeQ3S/vKi7IYTV8nkpMK+N7vgvdUwGgSlb7qWp2HbZblxHG4zj0XYTN8rSu3SDo0agBJ/
g2uAABzxxoUE964DbavgQkKUzZ/2xYPvHDMi57KpEFD3U6mhHyDK+GXjyIDN6DeiNgTeHvU1dzBj
2E4bGeFMXQ1jWfW3DJdDA14ZFm/14qmLTkvDcJTadL1qb1ATpVLFdt+PwYoIM1hk3EmOQEjNvrPB
f3ucKV9QOQFhIh93RajMx71wn1qWEpFjxxdWwV/0BwC1XGQUUklbe5B5Fq+e2C4j2GclZZVXzNlE
o5K7MRLDc+rkPjgzUQFqlfVL9IEh2ytkSz2KBtlFd1q4tYfQBhR5+TcIUj/yTjNYjOx0Sn/PWO8/
dbnZvjTWe4z7OHMwEiYiAhXddEcxSWS4rqKLP2J6lBzDDkaDqLip9o+2QN5J7gjWqYBG5I+5iynw
Gr43kUADe4ijiY4Uw6P09IYNGc5xir/dp/ilAP70c9oiUevvE4w0fE9BglrIV2xBwaywU3B0mml/
Rp+aX4++6v1SXAm8njAYx2R3rZFMshGp2k5YCTBX/BBua6JKUG+Fo/G1zH7WcSSsiwB+xR/Y8nct
jWlyQcGzSnPaXvUuUqd+tyryllzGa9RggUt7es/Gwbf/LwLjyNHUVfgKmtgHuqvRtXHgcZWt6MpE
8q52HS5TgtGcBsGmEe8NP0SL4tWzf9fVth2TuE6X5iz4xleL5E00x5eylRxtyMA9YZQcIP0PvQRA
aETMTIeWzyQB2g4h2sTSbV9wqSEol1Qpmo6//vfctmRKWhfJOBE/KhyEze4jxqzOURrp3HQIXhI+
lIfwWIHO2D66mQuf1tz7WR2sdGdpq5zFVe1NJMOCQ5cq1omaHAAD08RshE+inqUsejuQcqR174zW
/Bb7rfpERXg7femVjHYZKLB4tRzQiqwCwxdrISBp/8OZ4dDUBvU9FoBA6IwePE+uPuxGB3VssFuL
Qn8TXkPi8klWQB0HkvYUTq6PY/OKtrJrIw2fbIrTglvy0TyhJoOdsrw8Gx7GbVV2wdE3JNP2hC/E
sQ6Z9I2Ka24aK0neRA7PqquXQTza77i0lcAKUKi2Cm/sHBTSXp4KalmsgNxcFpLp+ldpeSM9I3Ue
CtJc6fdpOBNZ2065HqqCG40FPhJMZdgxB2CX+dzUmcd//M7SwhYgVKJKtEKZlvTC70zLlYP4kelt
4V67nTmY10wWJFLspkxr7d9CQTBvbhgwC4VzuksfU9sXWjQw+9SxqkftLtVfzp4TuIKGSWa1Y/e5
OvPi0B2yEqkI02w7bAR2HWY+w3fl39b81JUebD74B4LyaQNvHhWOxzkFvby66NLtTR8iSShEfcLg
Ji6dYmRWQDz4Ud78iheCJSOR4ak3SOPEZkrp4tppIAhZ+QSF4YX1nLavgkiw3D9Yp7UVlE+NKLU0
X3ci57HtdV/jjlBkA2NFzWhwCbXtLbXiTQTWfVOOTdbH4d6htElJ0XFNMTbJhJZIZdJFf9jSgE7/
IijCmb7BBafe3cpmJy76hlLZyuyH08CLet/kZ1ndzZrkL/ih/9BllUTa+FUmUEbA1R/hBviuYeKw
FlSXSo1QREnD9QuUymfiSjYeidvrcauaV0NqzpU0QqAhw2VYrTkA86aLPrMFud7Vd0Sma3cPu8dc
K8U2D7BERQFGlg0qJL8IU+CNmMlg9XU6xEGqz8MISLTuHDXr9fxfGAaa4r+R4g9Bsf+IPy5PIIMM
TtNxtlorD6oRxJMSK4JmA1IVfuXsW159JFCCwmz1o5LvIIAcgC+bWuyparzaMkfHoKA7s8WH02LD
5RqwNWsYnayWqoMwm02bDPVxIZX0CYFzbjB67G/TNlTGaODg/WbxSGkzy9qA3VmeI9Fb3qHCOPM7
WQsS4UxoTkCP+l8571QjVP5ym7yVLBs0VixAX+3ybDdXXsIs7WbpnAA5qbkgB8wGxZZYfByZSQH5
nOsR2FdMOecmURZ0oQbzdu0ktmId90f61oiyZGTF6iE5mfvnswGx31WHBsGLHS7X0DQX7UlkpM3T
pXGncKodyxKexPwU7jAwSfh9MNaMs4fSaBlAG2zviMcynptpq8Un78D9msUh6uLufUxIR7jzB3UW
sHXAqkoYvs3rKRz2LeTnea4mbXp9SAL5/YPBJflP25JOHAx4Ub67SAHVqdADuYkazb23T2lxxsNI
x6H81958zK1e4poaFWMsWslNKuFsTpb6cl0/wEG+LmIsqLObQbG20NsCJsRW2sLs7w98C018hL2y
RCBGc1rsii57/Is4YcsWkVC427xcCDRAB/3Nps9tbc08hczowIC/aBL31uGRfoxxu/s7+fBaFQo9
GLuxj91isEnYCtabYjByU/Fr2xO3dV4Mo+yxjMuvrgB97S8OvdntrarEukIhVkuhlanUMUrgmRf9
OCBoFoQ+y3jEjGFF0hyFE0UWELjsAwEKIj12W/oTYwNYsZzOMCCHqwzR0AULvi6CDz6bPu64i8AF
C4hVPBAGR2VIUDv5F1ZlIqXeMd57Aensn9GbSUL7IsqHbrT7TzM68nbUcpRwDkQe7bji8ifYcURM
XvRH0Ws6zgOx8AorYVC+uJtLTcKYqWHqCu6KrfT2lhzWBWO3EMlr2WsFUwMwuct0ZC2H0zXFQ6Qs
69sDrIL50m94VV/mNL0tAoUqcmBDYqyRCtJagMWO5dr5Jxw0AomeM9RFCnPZ7RpB9yzsAoMEthVH
rVGSVCAeftcO0DJJVgmfLPF8BU4tfliKhQRPnwaUsfTeDBcgyUm8iM5gsYIxsC7cSc2HRjy/gRuO
GGg6O4eSK2Ovprwz8DN9ZuejHkX/+Bqs8o5wWTbY4bfVWN67LaZNV4MlJatSn4Khi4YTqEwIP99t
hIgtdQbKJZ1gDzkvMlEKw7fyxd8L70/ZI5JIMLBe8s6STPAeafFJNWsGNt3jst9Cd/kUT9N5APkm
2kpask8IL1PD98Gq1JYZg8lryPtFM6TGmf1w953fbOG5ZQj5Rej0CNli0Arj3vgtmQMWwYECUMzC
qzB9vAsxfJPwRdKq+KAUDRxtbr2QniSMWddMf6g6AxBEty2LiBx9XfWbP1dAbSyhIz8w6CM/zA8s
jqyiS6r8XKNOpuCGoi3DdUMz7RRfFzdZMn7EGaXLBGwrZJTEUWGt0GcgnOSsAqlgY2uooLkel/AW
HS44OoU8DDB4qpzGp9m7UenPf8SFc52hBHRxmPxo5CbWIRdhC5nrb9vdbeDtsgyV13lFGPBaKhi+
7p2jt6CxeLODw6dA/dshqVLRCiBdYSN5CeCUxqT+s+MX4VHPtZ423tRTBj5w1KtY9Y5LTR2gWEKa
cCZbzfh+9Del4s44iLs1aPSFHAEvcsqPetYrygsE6Sp5JUiOS3ZJ8d4vPcpgBotXRjemPKatA/VA
1RlFftVIdnrfLkhIay0B2upAXs+fg6TMUwQ6p8QqeCPcq/B+pMv71lmiQqtjlU/RhYjqtt+7mHr1
mPUJKiIK8wGywYsfBcERw2Z5RxiPlPm+IwmUEAVq4ngr4fBI+68WSA08B6GzOyCwyHIE886iMHFu
2sTakusMLcq73As1ZzYeAohmTgdZ1sPiHTjJTGyqU2EJgTdadqzXWHqOKyOj1ReeOZmA1Pa3GH06
fuBLQb3ZHvOAvjZqo//rxd3YBCXFinLZiwrZhtg30vawg1eDz/k25qs4df3YuEiThAMbAzaSqgmy
sukWYIKnBaJOyU6BFWw3sB6VG5Knv5N3nEORAwuNcvnNu+LYld2vAxJidF4pMeGouh4sPOHbbifw
dczMnmeF0nFHIBqFfyiyRYTrPYJHU8XajGYvXKCd1ivbEB6pzCMo4yPUXWWbD6q9/Qi40i9fQwan
PmFGr22HGSEpiCkgj0cLUpqHak2FXxp9FhuA4GzvAKSLOBVOMfluS0aP4wNOOq4kZDqO03tF+poA
fvNYPg11cQrHDI29YYJQr5yxs8sz71uoWx9g2xHhN4DxBWcdDGbDBasuRbXxkVc6BYDZRYvrxIpo
xMu9COQU5KHUkCYJrfaDVyYObEabzAZBbrbzX8H06tHjazXEaZfWtaeix2wFZj5y1YavwTqJB0oY
hCx3LQJ1N+N9Uzn1S24VTHMQ9/esx7HTbTVuCO7qj7ISwOzPjIhYMBgux5xehcjKgUcZeWcGr9Hu
jKplYuIFeEY5qXp1S4WJzzC1s6g45KPjIaY2MFPyRnfNOSB0aGfhA6WacnrzK9lwwAKamnT6yN/O
Z5AVQ2sc5qi4qdb7Q9B/2ac9owOzaCpd2HwgxNkev4BFwAsNJLWMtwEZJE/ma8yNjp/UTHTyVShJ
t6W2ocmtOwztcfzX8HGmvlC49qZu1p0M/8WmmAFt3AjpmHpKrgxR2Ln8MO0JKZafWIhjlholw3qW
M5SMVSw8jNoKCFLrtu6LgoNfFuisfs/4xFYp8h2buVk7t0tQre0bI+4KkQt6nzDB8u2y5+rlU/4z
GQDCfJS5MEQpRlSSQ+UA/aTzRjt2pPQaw9eLjqeFL35mr7BUTgWZMtxeOrAIuYCQ/PI6nr9fW/W3
f7cXUJh7V1nrPAJFTelbJWvMHdlE81dNIZLykRelAPRYRf1pR7Z2wdF/w7k/7Bs+wFzHV3LcgwR0
7XVXwkJKvee4b45IHuU3D748bY61udMy91BHu+VClgnnkddpcNeHb2ZDD/tAPtQcMUqnuNo32YKp
/kd9olt+OtM16Lm1e9lYiCPNiBr7PpLq6BQbn0AEXDSYcLdjaffzIwLCLKofuCCRiN9NeTRsQpMU
jXxmVnVVtTbPJG5ApPn2rj14Nyh715bUEJihg6e1vY6fDdTo10MQQUL8yHWgL6rZe1X7fL2nAu4m
j8QwK/QO9Gii8GqAS+CrG5vZRP44jtLpba/XN2OZQ+hKRageoUZuiI0oBjBdRpzHGEQCzSCnnm5b
ZxZOMjtjHmw4ASwN5nRHXlb/jlezWxfKyxX0NMonP5Nm4ZbeDtoc2PmoLMApUC+JbUYC1ScHPDGy
JEj+zUDJvDGMOf2CzdCgUHGVeMbvAFBr8mBG9Q4a2ytISxWQvXSw4bwgiGSe5JBrgoIxhGCBDgFp
ZrAzaoZDaXKFBZdhFdOSOctwf6QpN6J9QBklCtSZWu6P0MJC2fTrspFChAQmEuWE7u9CXsHZDOWW
BrMlChFTHzqWQ0PtwvFfSnIDC3GSoTOS8aVFNo6KMqxWEzOnfMfAmUtKf/PyJrqYzciaReZeiIix
wtR1/2zUg+h7CbvvFw6KndxTI8XdQLpUue/4PvCsG1OFMgfTaQzP+mV008PKdl0gBKrEThSaB/kX
B4a2awJ/f2UHDf6RmsB8D9Yg6/wWJ//bGEGQB8uz4vEwQOoLG/PM71LaS8bh1mio4LVpOF0YtOXA
W6/KjooA3Mx2eMaweGRhp4FG9UoWLTuyoOlPEs7m7/F4O8TVR8oQ1V7GZl/fizzCVeRuaceS4AGY
UYChDylY/Iz4MU5+mP2Jo2PQbNETnmfjrXFqPoVSxpAc1ceXzmHVwrBRH2wGLh7GrHLJOuMgQX+2
wUDT6GeOdRh/J9XjiPZhjbL4TVU3vuFYsY/Say3oUERsWHGJFHDu8Lql99zzudZ2zGfqSREwEiV/
qMBiaWE1asyiGe0sufSVfb3qjLS9oI4IbD9QVParMt3UFw7EEiSxiapL0y0r+nbocQpPayHJRC7l
cyeUUJLQ6BZi6qE0qbyEUiZMjqxGS28f9Wbsho1UPJpDa/PPYArOQpVj+lXXtr4LB1NNczaZjHFK
iMAwp7vIhQM+6Yk5f0vQGItXwLFdk7rQxMGQ4zl82tuDBeRsDQ1sWTsX9gAvASbTpVFBXfd4T2hc
2/7vFGPAeqxi5zMh43Da5Ov/nsKd2xPatkNbqnNxVoYVP7vNd9EwU88O4SkJ0NUy37Mrm20PVMYg
dPtNHkPyZ2lOvIeP2xCDvRB7rAfRRYBHXHTsOdN/H5GIRMCVzHFLwBJVzibCUBm6Hi1htCDv0Cm2
PU3yPmtve91FGq5Mb2lCTnCMAhiyC3LJZcRlWolccHi3TkbCMSnl/r3TspBYpv2w1eQMfFfpp4s7
tCnxzYxVezPZy+tHalRuDBBmA0jUWsDbSc9AYtEtg7QwA/z5NvXyR7nFjBKkRW4y/GwH2OeF8ZCN
q9rwUn/yAvqk4oWsF2IikKnFgzSrvlV2N03+zFp6+oMcM8u4EUtM9RXHt+2ikuiaX3ZvjFwNNX+W
52DMDOiVD8fuEYaTMaTam6jD2D16lXUoy2fw3rQNpei1/J+Z8xZ+csheBJ981LdCMJjIdtas71QN
w82euRt+ZjHG+jC4FTOZJXfX2ruCiHE831E/5n5NsDUKFXfMoKxCRS5d/859Qt5ied/g/JGJolyE
78qoALpSNNuXSdfkA6bLxid1xL2bEOgX4ulmVwDBLyaVm74Y+wCMyCB9dQZd0gUjxsp0u2v+JWo4
QZBr78SgDBT1XDbtshZe8cBISMge/DXtLyMz7c+av9DAFGj1ppZuGQ6xpbjZkNyQeXgZGM+3PYy7
sny8rM4V33AnLf+7GP2xO5KOP2JF7VOMsaB2LJEx/A7GqWEDZrCwUkqJJWgsPfAmYdZC9I5dQEyy
aWeR6Wu3MOzTl3z8+/E+6NL/IsIsAJZCD38snVSkFsFFwmi8MxJMYfzycWl42jtmO2f9CAuTNpG9
xjW0i96QmzANaPnW1L1dV3nq8OxC9B7KEaxVkWrdnfNyFIFS9fTL+1z4zQuF8LhNKKgpE0TMK1n7
id6lGyADo9zWrdO6KXALqorGkVFYTWhA2KaFA8py3rZ32xcIt1nqWJ4iMxSv2/EM8XTARYe6brlj
daNNR7yvbbOQci/P3EZQemnau7YwXiJhcmGmIqbQ3QFi/rGwGRbTsWXOeKZbIBacj6xx5IK8BSph
Ly4205+4TQ22ijKZIJ2eHG1oHkiT2O9sq3y0J4MM/ziSnJaf33A7iMhsT7DXxrf1XrAJlkadDqjU
q1gGyaPCs13ESnsOE0N0PaSDA0xQYLFMI14TrqbJ/bM+ul7hh9KzEr+Lq/eb7YBDtNy5w1/HlfRL
3hn5PpKqPqGtoXN+UJnNpFWpXNEtECKE9E/tYIkGBfCOvUVHPBoHWqngsJSb4VS5LiEmz5bKSfn1
SZQVBmTCwJfElkTq/la5S05bm0jbtPnbEOU2SSE4OwiYgTmx4RBnIeLZ8Z5/ljm69jJzBqt6ab+a
8eEZdZ753pX0d4dLSpWVAeDgo7QUUPT4bgdufgqxz9UABzY4HyTpA0fyHa51Bgu1dkJmK/g3lW0S
ZlpdUYltc8V6IFJda5/RFc6DZTyNUQ7XpGOg3FosAHcX4I6TejKNMTv6l9hjKbj4m8GzUjR+v1vu
R6oyTrPP38Qafin2CdbG52mpcEqVSy/bSceW4WUNvU+VSg3ZC148T4FL83ku2K3R4vcgeOoxZtet
6MHJUXC6SZJg3D77RYenymz8TOxnaRux+oyqeWQtbdJBwKNLEn7A3U8JA5reO5vGF8rSI90tAEjB
64yAkTtyYXD9OyD/YVjkVkiDEmj9Jxcob/U4XWm0vPCC0mmvbP5vknQtXWSREO9mTWQqoWNgXuMe
EzTH0yxIayVmtu2DiffbUwaxrJI84lg4IBUT4QQcKriauOwhkv3AEvRHO82NpqPzv2gbB4YddTpx
Bv6/KYYO8uDPfJ0/kWQhmMH0uaHqGI8BmNFGbbuTpsC4r6ytdaY/Qq6Mc5sx5rf+VKzQuufMcbuE
yAfEIei/KQBnZzUhaiLUYz5AMhSzla7n82IEyvJZ1rcmf4ZTSgbryYV64dF27M/e7w48IuUIPj6R
eAxt6Axz67fK3V3IShhfdHH1Sy7/yNBDJuzUIOVd/wRz/eX+QwZvJ0GPJOcyB7CPxpPcktoMZl+h
agbQ6TpsCzW61h7lsbrnc3kXbJoag3P1rgv/Uo1EbzpNrGzcyTp+qK8dO0vdThLVaMMMIkO5maEE
yXZm6yBhq/rGMqiATAJ9vIg5DpVcbzVjlwaH8b0rXwQkC/IqAv1AXw3nsXGLARyPhQycIrO68ENO
ub+P85HPVAcbsD3OSGXMyxPQvA2vnoOZg5LhggilMrarB+LE9UbGiwd8qt1rBUHktKDEVGqAXZR/
r+d4ry3D0yyQxP91bzlQNZ0oFDY9Ap08hmBLo/8ZxIbtXnX2Cn/6ywQYPSANvilrc88Musm+Dwhb
e63sny0CvucMHgPak2ZqeaAKIuwNWJiZkh+SyrBinRN0VymiyhK7hluEHgZCBWflV/CTra4FMB+X
pqUmURh/M/RDXGvyUtVz3oPCD5oCnKkBQ3atb1sSLKFlz4nVsk+ikoSiOqy29wPR39EIBx2+URqV
YDQ12uX1hxGWptd/S1ee5mupFHFvv/uiDXnR4A6TkGStpms8C6y0O4t/O7FYsN8SdtirVbtFvW02
3As/hyXFFLGz8KcK0P6osTW117N1aQpkOsfhY0y6GwFjc+sU2cnPUktSemA0ozY0EDSR0SG69uh0
iki4kKZko3l7uelUb9ga4yTAdXn3kQKjRPNYOHjd8TkrsG4iGiwcnlYH1RCpwyk5deTBw2flvPXW
6zUdb9fHYeo/UrYRGw0/m8y1qCG0HMH71V2jFOj/ur3xoVmdnk6lZu/vB5cBBAXdH4RyqETKGqvx
R1S3O+E5pPbV9kW6eZCS5tRcHP72At0h8zWFcowacRi2ppfOC5bi2PT4PNlvr9mGx/LANTRjx/jN
0vgHPggKKfMXr71lAE/8ic6rfm5Y8H+eXXojOUtE368f1HX0q3LNKQL1nOs97zf9JGRtjs6Af1ce
TyISB2KXxSCSubry8rjO4i5f+aiS0RAXUv5uo3OyAVShuDlrQfze76vY+sq9GE/wIzmDnKBIRgnj
PPMbzCm5JySkdv5/dQs7H2GHGwFH+MHMAbf6eZSNn612q4hVG+WkdKm6/pchR7zuutf4FtWfe6S1
CjosA5AGUeUYQbfpiQmmpT6lw4BF70OEU1JAt3Zx6a/H977s3WUKpmZxZWwHjVB/06qzeT1pDxX8
1CGYKlNZiOErz2Wh5UXEj1HXM1Cuzi+MDplFUQFTu/mBVgU3h1JXcC+qFcokMR61LuF3HU76M2ci
FN5iyuu3tKkGw1Y0XWL3KWe3MrcKfNrN7j+HJv/sX3cNnQsD/VRbiUQsbfyn1fiZMVZKgSGCrZMD
gM73k6vfvooDOVFQsVcE8LERwHQ/BhYfOsWwpsrJsDctPPs0mIgSB1PXGn5UhWKvu2ZiQNL0SJVk
RoJR2NMMSh0z08O6EUprU87WQeL9S1rHcW0C6U6is1798A2Tyr9ICyfBGlnrrdgftb4NKV6KqwGe
xfNcWBlugSgj87oZmZ/Pdv9HAMJbIEd4YgMmgdSSXwzXk1D2NHlZhYp9do9+L43DlY+DeCMI8ORa
6AlOvDiUlOhqrZG+S/34nWFUh0sYMBNlIpTh89Y/pkZLmwyuQ49R9xB4GLEf2+bO6bqcrqSxcMf4
HAzze3zOvr230M4+NKl9Gk5Mj/uUzGrc8UCDFSP7Opgx3oxZO9Y4PKBFfzgx8CpTr3QaO46Hh/w1
fsSjTEJtLWdE6eWHhQ57cvZGmgMj7w40+hQemKW76j/KdaGP/qHeYhR0eAHscnEBG5Kosc5PA1IN
WjHEx8H3ghlUyFxqApRxFirxS9WUvbUxFFjlZJ28mNk+r+D7KQA/1aAaEamEWGR6POn08sQzm6Ry
AKAYitxImB9q0hENr5ZBuuzTWL+yglpx6s284wXiQCeJiKUbPsz2e7+cuhJAmTkLFxly7td8IIHU
5ibnG8eSstqHJkhns4hdpWhsQWdzvAqWR4Vj8SgHHGU7p2UUpTh+rzA1NfkiTKzwjg0WO0WI1ikl
s8Rqgs1eIetVkI3zbc8lHoJQcS4URqIRXssqbdCQpjJbcFHRGWfyw+WzpjDfb2xKlew6oDi8ueeD
RP/29RqJNmCI2ItdeI5ER8jiDwP03NuxGL5+CgYa8JXHUjc6Cpg+6K8cr5Xl//pj2QdwDk2QuCqe
ZffXDcarDOBqJwZn4Hgc6MwwJhmACJWqBHh+0EcqqT/Q/mYfpBVtcUqukXFxEcipOspJ9H5K9KVS
mCHHKGsMZN2eM0PSgeGNKsGvUjQ9kkehTdlhIVrMQkghcKdpC0+a5NQzEb7OhWIZIyLz3CcCvHHw
tdDf1j35gNZ8nBnYl06PjavXghkvj3fkNnwkE/n4Y3n0gyDrYIisJRiYH9iXtGk+XEyE20T3cOIM
LEWDJ28xjRVH0M+mU2zAjOnN1miECnLW3+x5kYjQvxsg2TZzjLI/fpHlTeuSqP+KT06Gamfac/2P
3+3qJTOfwTk2qzTrwlsZ9KNRkUj5C9QnxGO/z4f+Hg/eXnGV8hYaldaTjOHMZNZcreLetyGudwa4
NB2pmsLeX5Gy+fdy/jHctz1xLCUyyeNItjpbEfMDcD0GMgW1BJ1jR06DSL/pDWLDAdal4AIgFb5I
sMnsJzMdjkGpkBC9cVB2VuKERmidz7FU3CJq3BaYyvv4As/Skc2vlfDbGbEAh97e6Fiz48L9nXEr
kyMoNTlh+vCJTe9qaPaBFY6+/M5RwR3wkYpChALndtkBgzWxwOVF6nhUXQyjSyTfl9MtKriiOTO6
0l8AOES7kzmHLqXF3pftrgILMFlzhNZzkNAeip3IMrYxUOZQUUT+/jWv/QhBV+s8qbUElybO+rfh
I+n4aoXGED6fbNnXeoSKh6qH63mHYqCObV2hLN0ndYgzdeUUOiQhSstMk5h3xqQMNkJYNGBSphKS
w5ZphFNxnfXU7yhc+c/Kzk9Lq09cK5ejWE4A9ZFSi4yisIhvfy/DFLOUNaHVNLi5rWV1SVXri9OW
uCQKS1FMY67s6owZdO8R8JHXg5PIG3/SuWOAQY7MHs7Hv85Lrf/X5KAeLkWSC16tLFsf4fI9W/MH
LSigyN36v+0J+B2gWeMNj3teZyEZwsMNC44WBIGTNZ8y58mDspQOC/0s80g2wEK9fTS4bT0Tzviw
VUsPF1EauZ+qriw1ignpsGDakQrQpucWLCqHxL7qWbMCVJW4/fdSLTkee2kD3hb3xdytfepAjQ5M
BAm0dveCpIhf132lI1eyOGS4SMTXT+dOGpwxH5kH0BNbw1eQEeez3b0pXNcRR9ceSO+xwa7+CJT6
2DKfr9RVnm+xI22rtY9HzE7v3umsBh1D+2vll0/Me7f9vePu6SZQyE78OXqjFSYn2TaCIUscrLoR
gHI+uH/nxDlKBHcpoLatio1QHRzyT9wU7wDomOzqpX9i8qyUYhNM8R3C6h2HR9BTq9l+DrIWTQSp
cubodZv0Ei0OCbMVYVvTRL3z/P5ZYtT6m7NWh9DSQTgOBhnBiQ1LepgJqKh2hzYP6YdRzXM6GgGT
Hl7gt5Rn8w+BuFIQM1kZzsWOz/6a8Vs6bN9mtnZFNnzRaVnxziXEhoiFUcoKy56rSoy35lSvOrTD
G/Uh77zpScjBzcwyYmQpLX7LqhFDm0I6LtfX0hVjZqdEMXLH9BoSHAZuclYNfmwDUpLyXfYhXXxJ
jQ9yx42H1YTjZtVdRgl4W9U7JCWA+0PAT/6pRZEp1mbXuUKb/0NrzAx2ZmgeaU9Bewx66UG1xJqg
cY5Tm5tukJc/T4V1ME7L8/LYYSXKHQc7xEktfywCOBGxMo31TAgfs/g7QyZocVAOdhtIqEeEFgJu
ZjP7XnBYk4iaATtkayzZaERARWwMWTLtPh45FCjPAVeO9cz/clsAt4DeSzL5SL1OV2SvZqIVElGd
E2JIiQzgLTW4TV0161Reb6uGcEpaZbWLrOVduwPO57mOBzd2bSOtWCEMb3zAOACQfRviAo/GIlTw
bcPuK8ZjptlL4SrG6EBDJD8JxM+6ZkJEodTnzOU3UyI6n1/dTGRpmdOg/UgI8gqemqGnms/H4wkB
uQHFM6NpN4mFyEH8PZG7fbXngA4nYJ4tfZF5l2BXZUHye8C2qbGesynf4ZjNCLCp6YwwpVJhT1le
KiMHNxIRNl/zGtJ4YGOZKxD3UyiA8l/oox3Q+DKk96tBQ80OGd2CtQwY8d0XLJGo+0wz08BOHr+K
FtqAOiM15NhE1a9qP7RntyvhO1RfJ/iUWDe6gSjh8uLzMlGhnGpkbY8xRa9pJGBL2zjIk8HgRuKo
F0ukNcWwnohs1ZsYl7r52qjGnGb4wNSHNQTnSMVK0XFjFr4ZmF1MlFQkJfUKNt97SahehgAmFOVP
Y7pZ8hS9Tt3tFrgca0XhcKINuljla+ooZQJ/44RwFa0OW+RQsUg4mn3W89NlHhjR1mgpz3Qx4k5L
YoA9IkVV6h5h51rqbAwsrYYl/z8YZGvj+J1ETIKBg7m0eAhmkIFURCiGnW26pJnegplDH754X0X7
4xHqGWMBpZ3b8vp6hXKiASH0CK5MmjFV7Y1P5yRygcdmZtaDCrCWiWFRRQ7avdnmkxF5Bd3CCntY
mvb0dpSGAf/+R5l4s5CQ4+6zlPkSVHCgp7Z/BFGiLzDH2GVz7Jvmxdq7KoyuLX6Dr/eXZZQucJXy
a0vFAaD+5klOxP16/5Axa07oxShXha2KWYU8PtIaXhPN/8goJ4vkVDH+HpZqNdj158hHKakIlkmt
K66MfClhb4ZEr2LTIRD0u65pN3L409eTXPDc7m/5uklGJR4cBRRgUCe3ZfiKWDu3QQn78YtiNbKn
bsJ1m1KWnyDVw720X2TykNZmALZvPh6pVVvmlFhD60uGdUS3pomnicQsuPUdAS1C3P18aTQWRdJ2
2AydaqVRZU8XwrohVAtUpx3sVk556wush6rLKhKMMCgzgISCqg11QEdQGGVHjhVL0NwNqR8xDTAr
c9buP8FFkZVEaYTcwNybS0lH2tdxDc4Ac1Ni+VpDLseod/W9Hi11teiXScIHKu2NfywiT8DumgAw
/SsTYy/GIs4w2jvJqUjP5ReRg2JUYrMK/YuSn4JvvoXP798lPP2JIidBl8JqdQScNsp9x4eSkpsa
2++CNkGy4I5uvhK4OPwP+ebO8I7Kdb6kW/YZ1mAvJ4LBPKfwt3/l9ODi04n8YbvfiAneXndOnRKR
thyIdB8hRlc+rLY/1fd50BSapZzdn+8+8jXF2TqZxq3mj7olqAusesS1s+K5VN3ho9RGbLC9Wvj/
83C7b8b2K3w6GY9nW0v14iGkORp6wUwCNQXzHV5ncM2dv2uCi0BtWFfM69rT7sTDhj80/gJxQ5NQ
Nd7FEOgGYL0VrNNsirieTf+GHtHWa5EXyUfiCLurCztK246cpzQR+xDJRV3fLnbBgjy2nzkHzs+c
JBoBRcnUy6H1GMKUH1PeH9mkVR1zkOU9kPHzL5kHyaf6XpHQo0pImbcHrIcmSb1WTt198Od+QUJQ
mSaKSCzhxJ3TQ6o2XoynUZcPYAvUM8RauDqFtO3SP5tU2WfN0Xc+xMaWZphtevldpEbZDENJ2WWg
iEmQtO+HDOtUJ/6J3vCw+DjsYihbvX64z+lbR01sa5ENB8eyRYfdqujwjFTrnqi4XsPDPwS/69Am
7in+9nrK9aVnFPCEH2Pn0rVDaNljoC+Nv2NVsYaS0kGkA0WAYvUu1ItqRS60XH9AL0aG0KynxnWJ
6U4GAU3ymvmrTsQzdXakLC/zr+dkGnjshvzLGtbFVY1a7svk6/maNiqK+81WQ+8AEOAducYzQ4wI
9RVynni6+BcT1Z4BcOOhKHIaVSkqJqG7dLKiRAkx2Vlie3zp5ehHY4QyXQ9Bt+gAg54KDeGjc70r
K8/z7Yvvcwv88h3tJDN0um4uXqeu6mBZtxemxeVve1MnvJGfuCdC0tq+edXCjH6c5Ck+KeYKiMMm
0kw7pJl8LQWa0A4A/OwZVLGrbLVPNhbZyCePzRnVtbHYDuYigvRXwiTc9EzQlzA+WD4myett4kvC
beDPo/pCVI+fX5w+izcBj37Qs/kYg0UfPVPtNHe0qBfSOaClNuyj/B3V/6Ld4eSYTOBdwtkoO44O
mYGri5BeDkFkEHZrvz0uySctZkpkh/bi19pJHcX2rWAIv3/mebNRR3M4Lqi/BwlyqujDGBgGTAYR
TEXFs3tru0107qLCo5705noqRBVZE0zvTlakW5OLqoV9iY5gy+omlAc0JivKBpCIuSlD5YdPSl11
aFA+QfW7jvBE5XnOOlTgKYKp9L8nRELnK3HrTGrqX/fGuToJcUchKjQLJKnkfO0Cn5tUNV84Jm9U
voBvjayRsjuVIrHXNZKhOcQk1q4BwngvCSOapA7tQyNNwZ7ZruvUEvBONr18I0tm2VzVX9YM60DQ
2sAnlHGfBIwNoMSt3asBTPAQNPX3208gKtEbJuYi3BlVx9okpicQte7KPZf2N7hTiml62os7nJVk
IL9mZc2ogk7wh+4blHzTqUB4b/KyBlY50FGnNqil+GCsaPJamEnTBA7PXUmq4egU5e4kTehfHJNw
tswYQStXsCpqA8Frrge6u7duxlqXVSCtlmTnryQLCO9vGTFwfShQX0UxV7qzPS2LvgA31gwRZGxF
V0+EXDwu3WIpkK9cI4CF0B2sYf1E+D4+dxRBDa6bc29ZDAFjqiASbbP7I3BJbLxzMcubNmJPALIP
N9IJCafJgewf0+2lmT4ogEgoI6nBSFYKqelKJIaIsFBz4qMT/EoUfKtBb+XtTXQWFXzH//Zx8w53
6GgILEGYi5JHlNkxBWC9sPjL4l9EZknT+jhcyQdWLiWuiVP+lh9fcAPWUAWy5qowYdJIeLRrjT02
QEh7BDfr6YZ0CQ9gyeGr+xzYqQ6IYcnGPFJy06a9ZJFf6/fJhWbplLTFmIzk9hFgxZY7grtwDt5y
5rdMsDJVrAidAXUz8xAOQo362Mk5J30KNDsDePHR1Wpr73Q9FgogDP/jEsTwdHQxK9Pu9+aPu2ha
G6ehsBJq/PVgY4dHDKDoOcg9pOZDqbe8u+eaNmVTjI6ySmaP61JJzx38LuXEDwoEWWWH54en3dkD
rRviedjxONQAFrkCANe9QFt1KKGY7HEXLAor81Lijai8pE2aLyHgSCYARP1oipgj6tdxVdNt/jtD
AZnIcncxMJGPmQSRIcs1JgqJafwg5K1TKiaL0C4BobwfXQv949GWhCBwwb7jWTB+qL2JBkhiHKAP
OVrqtoPwi9OwNcdbhoWZpdZFBrlbjmhLwmhWZag18kww/H0DbvOgKI9V5cBbzlVQDe/qgB3XM4f1
ztJsU5LRf9uU33L9oX7MZXsp4mpXTGZIqwkoUXrekJJrp6UGVeDwEyMkczMcos2LCD55xgJCfZWN
zHU4bD3N5Xl53IxhyrENsWnIk+8dUAurIdctULaL/7VRMU1yQbpbqvUEwe0zb/Vsux8EzLE1qmO+
lR795uGH8BpEniA8LH2k1A244QoZCyPzkVSr6zUY9szhn9iyY1aLoQVIqiTkx1tYt0m9li/qjXDY
D4lqqmirHx/0d+VFbY2wGqx3Cczb7vPLk1ZdZ3rqxcbrh6t0W3KGWEmsP6/KS0KwtlqOSVgTzMzO
del/cm2oJ1YOH8xtRoerJxvfEbYdpPc2IhWca65z4peBpbou5v8j89Vjf4+J4qwtMluiBeMDU6U5
coU2TpRUV5kqzfQammHJL5qjZAh1St/WIcZuJyFddwfWhwaw3lU4X+EqcnH6sL09JNq3gKmwm9/q
cgASb5stGzgl4+SjZXOEP4PH5u2DtWTOI2eB+KPnM/6dC3CIxpyzPEwsNZ9n6gOVdZx1zscOCMnb
M1Ez09ZdZozv4DVMDnoXaOMAeIfah3BfxPR1KoVZwrnUC0amUB85R21dXVr28LKlCntS32xyUVLy
t3QRk00OnawAFuUuKMmxeVFNTQGuJG55oFLAM5pQDxrqtH6DS10DU8gZC6xUEtI1TbPXfxCM88BR
sgGvX86ivMFtImNdKdVzaLc0RL0dTKys7P/rQowqz0pYO6rzm8jTe904W/6pBG1gBE+IPerYNJXH
EnSFQTr0vfEjXoynf2aD2DojCv4j3h3B9Sbw65wftD0xdCEK+ZD9Mbqa2eLRBsAMWxkbENhrkUkd
VsPmz2TJXQJPvMxAvYMAy6M9afjjyX8lGbA3Imfyb1ym+p/zYl32Z7wKhEU2oRi5DCNujOWM98/x
aTpWOZ3V6unMvAwyMBtLy7FsusWxVNiUsbZNlq0kSgXG3IHaZGRPUOOdCs+ZMzUOhDtkeiT3My3u
Zv7I9mCdGG1ckzi0ObIQZekH1dRsx9W9QO7GwP7e24vuSWWsyBkLl66ioke601XAc+3Uh2OJBL9e
zCFJs65uoZtgX09EveSlmjxBarpUGbxOoBQULQ8Qk0xLGbJSB8XDI9C8gYomri/Ctpexw2EPu/89
xOX5n+NLlZdmI/XvlcJ1xAeWZs3ju0C3wockQ0TLxSlzia6PiIJSCgIxdVzoKvde4rcisjMvbaBG
wJc8VXIwpTkoeTfCk1fcuDCFHPvdCPEdhCYPRsK6pt1UfZIcCzSPwLouftznmOeKiQDf9oNWU3lW
kOCme/b4WcrNde9jjWGfhlizTh6iXmlNM5sSpNKrYkAdLthu5Li/+1F10NJg0pGWOyEvpPUIpK3n
FvRIhqJ0X8hj6vvBpqXUcTyA3nwl98K7LpbWRhkCOUoQXS4sq1V1a/e0xcGDkByxOtU4miYwlNnu
DKuNIIlrZzqMYJu9CPys5Jp31zu//9z/6363pKjhcUkbUH/wQwtInVFXyL/BD+Iq6KMz365SvEhK
v0ltREIjFX/NJ3Vn3oAYc0d+GXcbnqzz9U0Z73dg0KC3ZMOlwGx0qwCrdLJKT+xsjx2km5K+Y7Y7
cUf1XjhTspz3T9rW6RAQLh/rBd8gRZ39wz4q/0YEa4olZ0a4uch/F0tkdIoSZWtH4uDlYBnZzoWH
SMtC+Er2VIftMVpJtNBqhbULEmKxCTNBPppJIyVALjdHU9KC8JO3QkvcoMOEZGOYdlgKbPegZLrI
44hnYKELcPdIwxBVgYiZ69R4LytXl4WK7v9MBgTmfBzQsgP64yBRpM2B729rnK6al8ObxPcLqewO
BKB8dGXdhiyR9dfM6Mtx5+I/pA6iXdXucyXzFrZX+8PeQdIIteXkX/jC4DfOazaSPyIQNfPW70u+
cmwQZjEgGlP/4vpE91SSrxJX6sCsP3yv/wbmHMzL13yWDYbuGONpZIWx5954tIHIZI/drGnAAcRr
WkFo70HFQaO3mtQIA3e+WjASbYaA2vYWP5Em5t956ukzO5cgn5BFaZxhOBrYbuujZJhzuVQ4SWsj
m6R4Csqu+k0MlhnNMGgQXNWc4p6hw85pKUEwgEK9+2tIW4kOzZsajffR2HXr8w2ZyRa+hnVGF0ZB
i0rYANTsIGfrGAhozjkNXmi0hoYNmEaE0r33j7mhIxq3NvfaTftMqqOBvvC0IvibDdp6oIjxqGlK
zibOCNigPeauxJhWvQIR52o6SGFrjSmxlzN4TsA+yrfhZ+0s+TBHTmk4JIDytk1k/+HVikX+rVFo
uNz9NRuTaEHKsmc95E8lN7xtQ1RRIaxNACZ61aObuo+NM2Oj1UNTvXwd53Q/xXRfuO7eXrXmZJrd
qekgJSIu7thlCTuDTa4FeWB2Cedz8WCXREn1tVYFTHbryhiNhzKxAja+uBg5uOBXGoiy22axM9lg
ns0d3MdW+phdcwrjws3FeZnN/QfiOZOu+F/QWOb7gTiIndhefDacx7eJEIDI3svljL91NQCU1JEj
/Ya2Uh2fUAcQ30wG1RrvMtZo9sBckWMLcp9Gq99ijc3yHjau/6aOEIV3z7Fiq39zN4SqD7O7dirW
mSCUkkr/tRYttoUbUEY2kQaU6FirJ22eFW0vHYFwZD+7zUw7yCAhteXGtokmarAbCJroLitm8f0B
UifSOC8jAZotrDwsNhe8icDdofkEfNQbCw7bFpV/VyAuL7NLTGzUjAYBh0Oej0IjzrVJyxac9tWo
CVJX3FcIp4dSi/GVIu0SD5QuzbfUWT+ma+kixsuOCo7DLLr9Lv58COxhl0y2FXds79Cg1PlTPzXi
MnjAkp1nDc5Iv6xYWkgoWhI/qqfqlXKiCA7EdEXvXiYw9cWOdSbqGKFzF58ymIYo9PeXMFj33kyB
90CVDXiCmUSKp64oItacgPbZpy//X/b4XtMWR/8SF9dt+qM3HjNdl6ipTenoomixF58sTjntvrXp
lLJa4N7P843cw0ALdjDe+YN2QRHel4YvSzAnm002Qqbhfg5ZOTCkTPf5S4xO1CgnjnY+SpbePAvB
tHGt6dw4udW9JINcsSYaw7P5Gir995xdqyIuRJ59+U/vpJiCB26pTEH145MctrHxiI++HhdAB/s/
/inj/COTWZYvW3qbYjiB95q8XwplbUZFl0VZQmqTUZLstUQl0cQkirjXPoNStC4Pd37u9FnMp/+7
siwg1UiaH9w9sd3HgVHr0bXQkajQ+NP5YIH+a7wJdsfb2Hg2plNfw4sIQYaJfjLjquUSbFJIzGkH
yP78PcSQBpEMmzJR/xHF2pGMGUtZamhPMTp6NURBhodT+Pm0MBwQAW0mU2wAm9Psr60Yc4NMxxoA
HIlBLXrXA3O7Uzx96+/NRGc8Be7zNzSqo9RjsHlI3tvh6sysLKWFyB8iwpyRJmRU7cafZDjqyjOG
2Y3UC6qJYKDM4vPbuOncAmjCmkYLRVXhIOyICP7P6uWdyk8+3OqJFjFMQp2cobQbwb7E13MvGfss
awphDLHxeapMHFNGpc7WRLqB7MIxhBMHYeVb+tX8zkHnP7efVGRQe09oqGfx15NWnvgkRwHlMqqZ
wnE46mThdAL5SifT8WhhbpCbU8obnvDvtTM42+Q6VhKs4U0Qz1bcsv/dTFewsJqdCZgo23mW/aED
beZ45N7GYjSSJXOrO0Z6ddWyY4GOrStJAfX2tLRrFxTJPmzNF360WwvZpXOzhK8KxGQG+9M/DQvf
8yvQzfmxCG6qFdPpIZ24AYXonCJTzNxN17twMaJxaF96kAX0wLKG/k/GFZWVtycsZX4pumSDP7Cg
9YFhhxY5EzNpwufn0rB6vNUuvk+f0weiC1Js2RN9f6RngsB83X00Wnyah0xoOqnMJZmFUlwJu1f+
yDxWaI/XORjz7WujppnjTSb5FZpqcQ1z63Yvt3chL1yI8onGuFF4XnWFPGBJ70OALgVIlxiLNHLZ
wSKnXLtABn/8unOPj6HO9FMpnhOSUo3GZu6cm/c9gJS/LrbvZ4/SGkoE9imP74NcICpvy4o0KzVK
2sYs1zk1k2eRKbPGYLBQMFiZ3jBMDxr4ngbZZry2rKZfcUMoPYfl07DRz3iUim8Yq+D0z0DUMz0p
/a97Vp3mQR1VIK7RaOqmViNIaG+41Jyh9ztPhlE9mEMcXuQdibPWEqXG7mPsE1vgDjVZyYzOMjeg
5cwd4mLPuuYy28SkVeYSxSmNQnNC43yb40l457uswX3In4hbkD5w8S6rMAmF6UH6L0OikefzTU+q
duvdzby0IKiFCYZHZOrwSN6997zLCJwTx0CNyiTSuJGN62MbRFT1+mZlUJToRfVGe+Aa5XAkHrmP
FfJpGuZLkWougeFFaT9ww5vBdrRBC2pWwnuPsz9WYqNhcgqtmu9pYsvPMaQTgc/A2RgyJLOQ3Qat
0iyVc2wf59W3CxLAqG7mVyq5ABtY/fYUcy+Yu09b0kWuYlKAOQKPlSWEzvNOPpx9VX9DSCsf0I6M
Mciucu6iG9br5S4LrD5R1Cg9BMPraOfDCwwKQdHUmjnwP5Ohvf2BoAAlZ7OAW0AdTFkZxZO+j961
vn1/vOJ+QR+F45V8kFN/3PIjtO/N94R8ZT4U793TNVkYNJuv06waWl7ALCfiQJQprUgiazUPpK6A
IXa0v81+nsgpdmDpLv33vhPsYCAF+rL31Vm31L9E6G+RjE0MaCDiknM4tQLLoU5sz6/XsvOnN07g
iIgqtmBsDiDKGdb5lGx3D3toVO72WtTP/nXycoc4GrZZpFNSp/Y2KNLkhnpmrm9T5BpQlSofX83h
gPUOmBE+3DDe5d8UqL7Ur62tqyuy99EOckyLHy01jggZoH0qeznp54eFYzQYG/2BsrR5bgG4ojyA
JAJaNnlGQdBldiEYY8kAlq5aVOcv9ZMc9Uir1iQfNz960jZEJeYHaooJYcJePqSxQBz2LD3piExv
MvmGGRrD6y9hmAWoHh03whHQwNCsiHgrUCamOkiW/03fxIlGw41f8XQcYL1mm1AARuM7dbgkqV5x
ndnQFqoBGtz8Se4f7LBuiuDusRWNyrbHZWHaNTDhq5aa/PGkxqSpOPCwJ96eHs780FaAmUItQQI3
4uDJb1PrU+MejkHQaawvPsmAgx8270zw86MBEg2Kgs5ZKmB6oBgXUL9MYsdLh5tIFOpET96wxpWB
qbIZdhtDgNgI0LayFvUgEBPAyNg1pKfzR93+DFPIchhGdA6azb4Zmd4JB6AxmS1nrPMO9AAuyvL5
EfjKIAMtktE6ChdhKnHEExPELILHCzDs5F3iinWI8MkI4JzAvrzoQRjhyCuAfv/Eu8yiIbVryXlQ
TpTz4XUeLeauc8Hpmc/6RbUPc1FK7xn4deTPgHr2xAlravQmYNwObYujLsCEvp0J2RYX45gzCJCo
0fslmiRkwPMSlafQmsqcYfh8EzSbdfZz8k7nI1Mnycfud2k7KklHPlRk4/F3iPnxlHb6z+2FewTG
+m5wLMBeu80oXTQj35wZzA9FpjzCuiW5CCbbtpydswIlanmRBqirjf+tMXSZVqLrpie8V/irhGsr
UcYekscNKPQgO3AqEAKbJHuqBaizT5jMx9eDQ7H0TDbsgvS+6rN8fsjkTQO5mUvqLdwjSv+ufQ8F
Z5T1Jc1AFH7MLlQuMOm1sh6nNtsovCEjB632OyXD3MoZwbGLvOi7acAczpS801vExQkvPW9bnDQh
vJzWfNP60Z8juS6P4ZgYIl1pgRjsoJUpwWyjOi/f2i/1r0uMD8MYFGRAxSjOQXv2weacblKpmAFa
zBFJc2HuhIdYMyIK8TBa2ZTWMXm6hPRI/F96x1xDviFxm+gS7s71hyHZw9ohfsf9bo/BKzr/kCAo
jUY5LcVEOmedmul6SdvBzPO3EJPgjdqJHL2rGBVrlVrLdsSuMWPkJRzc0Sl71AjOfNxRQnGF4mSO
+jjC0Xm7xXPlEK7Fe9NVbXe7XeZYWCng6jdWuI5DdgYHpY1gU0xsuO79+jmd31ngn5QBSc/m9rd4
0REtPRYJt0VlZSLQgKReQP7huzll4g1vPEnYuzK4ZZ7OYsWC0fYXAU1gd5tUGQw2qL35n+I2sbPJ
gwI1/0delmT2Kwr+qVL9jXJCwDoRJu1wnOnfIY0sv54POaOfDn9/Hmb8523LD1GaZXzKGO5Jukq6
GtmVLEmR1UCk8e42FXZ8zOV4JQMZzih+6k2TmdrXJiiGGz/NPxq3kWmE9cWEYTpQG/B6RXy/3z86
2zcH1NT0geJF5P498TAqRJLCKtjt8sE8JjCoN4TDpVKWOkkoYKKE6CoZbHT+//GMrvHb9a6KpQ7V
KpYOmF/aOuvKwKkpTeN8RRV/FM5dYg8NIF3B2900yP2a+Bgs85AttKRk9H0ATFbs8d+JcvwGknbt
GWNupo5/csnmUdVa0vcNqLSvreiUKRCe8gBozptiQm8hogkJVNIObL7VvgYZtPVMERinyMlwrHcY
RYFeebhNcTHJW9mLZ1PqlrLna6jk3f87x5OIE2V4m086hbLnxazuzRDZ7KeKVAJ89HX1brOGl5u0
MsjJq5dyfeGrIQVbFWJxVrHG6OteISfbrWK2V7O0HTmtIxMqIGEenlLz+ntlmNh548r2Iy0SOUea
+uS1UwFPTDwyJX/p6k6eU1RAgP6v3yK6hn9gOu82E6H+9xdmGwTR1Umi6vUXYK+cd7iai+pyMdXA
kyXo0WhPeFhvrfGKfhuOMnaNZruDHvDBj/JPlRi+ScZy4dKkuLTyQQejXctpUExnCJ+folxAPuAy
ZKxfS46dkkpnnnFqOxjWO5TZzDEbElhIU8OUhIv8ktQk3ybktshN2JWIA8rshkjNeS3bKvOlgd77
0ROGAk9U+AUHJtyrVU84FHSyJa16lnAGZzhiSfxHVp+1hKsmoVQZ6V/80QlU+QOy2zfFGHqULXLA
ivqEABgwWEsryoYcfwil8ByucPuqE4Nv48eNagDLP4SGYfoShjHYPItaoJ9b5C5nyVgWTKyxTt9w
gM5iejYLVyjHzoXYAkcBgNwAnLHp80s9fvNW2Kn0nSh9flnF9NwP5oHRiRAdfGV5o9hu/y0B4e0G
lm7niKpNXpr0mMyGdDdnG2iPRPbEKPeYweoKF5oxh8g73XalFEhCSB+kV4aD2HZ8Io1eQHTQWKk7
x7Y3B+nCNZ1qauF9CpyadhKX+DGqzFjbPW2X1xvvUiBSlMpEb1imaY+oLIiQQ7nYTH9VTFRJzz8I
93S6ylbUhkHM0kA1pQr8Lo8i85MheOUUpeRAsMuo0FeFr6SVmZlsQ4xMItvGw4YGmayDr/mAEvJc
8lAWd3cauVa0csCqo/2qeDzU7Knmv3KQbKu5jtiF5eNpowSDgS95zZYTFkjErIAXLYfnLEtdkadP
ZEEMhs/JvFcQz69eEehorneSGw5yEFC0v5omIkeFi1t1Tbm9NYhZWVEk3szHgZ6wYi86ubbpXGTr
9K0jVBw5ZfY7wt7Gabx9Mr1pN0z+zCE86kB0OLw9d5gIkDNE5Ph9XNY0S7Ss1CfdT8Yxu+Qgkj27
mahp2ZAn8aXxKBhS1sPm6Uv8brwE+fdBtOr8bRrRjzcAOuGMZzEfE/hKJHkbL0uS7iY1tYapMMXp
6F4Bk3KqJFto65JSyDUmuJgOo0sgb1C65eCX7rMxb+mMV+b137Z/Q+2q1W+nqYbPY0zY14vOBe10
432/E3ezDvyhbMoZVJYVdiIwK/eF46Qvzuv6ejEX5ELb5ni9FUjZHa1uPa8r5v7Wu4G7C/MM/Hhj
Goo3Vo1R5ZLSBmLM3X1xq6IVI4GeAPfPM+2fGvDttL0Xeqq+SogWtl1EgWnz5HMlkLwpsW672rOG
kpWK/CQN6SPe1k/IdtPCo6eFBQsrftzv86WXQjWRNkWcUPOd6BlpAoV5WovkJq3rCFTFBqFrSLMt
v2De5hOt3BzRLyj/YuT5iLyOv4H4PVuVZwDMv7kLItwznaTVmqnYKVuuv8hDc8C0BNxdBuh9I3ac
F/btx62O2l8ua3L6zuuDs+B4JZ+L3aWZy+/iOatZAP1+YD62ZgNxWsBqw2gl89l21Ca289yaJwzp
63o3eUYWgkJ7qxeCbPzpY1bTTh9fq4PIyu2I/9hUCAdDRB6a+5SVG1bcPOilrbbRFCPXn6r/RYQu
2lH8WMIwgUe2QTU0JtXpPZrjL/jecUmBwo9DVF8ZOfw96SGnW5wCrdJI+vIA3Jayv0P+TstIYRQk
xakrXAUXTk5/CUHY7IIIqKO/p3MoXtaVf1AhAZ5z8riFJrap3qT7NhLd7B23JNSSil/vonwDC+M1
wnrYcVXAFDWe+CbLo96T4tM/GiERHu1gtjmPyosoe64w1IZrShzEnL6DWRz009boMK0n2lL6jMN5
kLLdi+JqGrMQumraOEcyoiunuD2PVVCxRrcSa0BkZ778fkdzpsuVACr8vAV9hxmHt/ZZRAD/8zqv
m798RQMJiuXgYSI/GHK+nhheyaF6DENFCeb+f/a+qoiDSLMg9qKIS7l+mJdUge87kBi+QCIttlDX
t2xhc1zqZbS0oii9VhwWbL3c6zYiDuZbdzl0+5BPBbKOg/AE/lkCDG31lXJQtiiZQrJiRUgikfuQ
DaNPbXRLZwPCR+KV+Utjx3TgEB38ICl+21Rku3i67FoQ93bei0AJjCHzjBHRq1LnYbifn0n0A7At
i4CCG0OJDlYRpU/sQJpTdsgkyU3UKNbqOZ0P1zOIlZRgHufQaE/sJMMsC4S0mUPaB2W2LdJc8I46
7lQsTIzOM3qSBQxQYk1B4AzGg8FYy7lwi8LQGYr7O8hLWXb9MzSyLM7be2rxRwRyrCU8DJ2Fi7Ht
/kwfOpmM5N72v2Idmb0171Xfuhy46YgJtMKvJ4+fkpviaQmdIFsTbyxt6mM0W2CJM2OtK6nuegSo
4EGA+hrSQMdR5u3I4MYu+pSfWXWTh6zEAzvq9kGEyvorWOrxkUNlu57jSH3ziKHcBK43P9fMLDj1
+wKmdTtkiXOxFWamw4lCxUF+orserJoreWzEj/Cheptih53gfnOybnp14dxGV9fVso/1nOmy8/55
XxZBCtI3edBZyboSNJAUoht93AcZb0TJu4lUZlhNAU7DG4nPMolq3bsE/nSfENLdi+SIr4bC2BF2
fIniYnZkK1AZiDnzcvMvEt2p3WNuFq9pazLSnT/Jpoo1iziiUpxuPfc0/j+ga41rcQkD69lh9o78
5lISsKi4vXU0bS6UBj1CWhOe1Qabar9b51V1gCH5H+9VJeL1sucIKO0XKd29VNF9XZHm9bb15fMx
nDIOrT44rSjodSv/X3ykLIkqxv4rKA47/YcjO7VuuyR1BEtJGC8Bnt5ktPBtU8bS4D2Ukkofej3A
z07+VBiZGC2NELM/bQ5ZGsu0eoOUegAk2mBNaBvkUIacZojen19LZo64ZCULgdEgGCeOjtQUTXFq
R876c4Z4kHu9feZm4i/yFgXBRSmdeLLwnXNlvkwx1Sqycqa68cI39r5wbN93DpKA7ZOti1toQ3fj
byHDBcwBYMQ415Eah44/sWiHxSLBap0P6Uif5brwYbJpJBmnNeYRbOFf9AhhavB37b2SQj1hsiM5
Q5JiKxGQxgGjPtbQCUqTyZ+WpCbWUPmUeVLMniVXpE/dCIxcmTRgbxBl+gpGEqFp+htoFsAYIEv5
ehO0b3pqaYJ5L4HUkuIF+8j7tPAyBWpYMj7Th7n3r/ye6GMJZrE2AKvQ/4K6jEqkJxF53J9CgxAz
xwzknxe1TCeL6YgS2CjbG0rcByKhUzXpAAr5L36/Nu8Q4FPwNsk7SSBdAQGTdKKJoFGG7LyZsats
xFX8jiKNlrPS15Cdp3RZqDopZDoIYm8KVH66g6mcpZmU0l4zy2utsexMgAbafY6/hhhsb3jzFf8b
G95JaYvhPRZ5D8U5zmqBBW8biln0oVndOBAhiUJLNAVx1XdR7Rthb74sn+AoTzV/B5v9HMJuIP4S
OjQRC8ITxzAPJP230jha67IBTEJq+nTAQw55BKdlF7bW3DjDQLCaELR2SjNgM0qGvGfY1HBH3Ycd
xN8kwjYIdv46/cubKiqbFRyxPSlqtwzD4WRBTKd0J/l3C9qybmlo1vrgAZmaUBczZNDK//Uki89H
XqWN2/zr+Zt5LoIB2h6znwgx1C/eo6IHvnLMV2x9Gk3JOtYH4t1BleRSOb38dDpOihfTp1H5huhq
t+V3ZmtzovXjpSFpyBfkuVfhKmTQxe617+eKvGFN0pjPROetdn1k1ecDkUb2GtVQ7KFO45LXuIWm
/7i9lWGgZkA7IRw64Le6DHhrQ/LOaJTW8+4tSmlGHNces7Ip/oUTBxQ2Xsihs863XTYDTGU5iPs7
UT4BuJbiss6PeG7SC10ilBqFx1m7gNeMz0qVPLlXQqEdSATQS75JV3cobYZPH2EkMAo4bZ3UfHtq
UC4bzxZ8rhngn7xgNRRvZH/cgRKDc6FRk+tus/9T6dGOlDW5hjijvjvkuBzetjCR3ztFx33jpfgW
GipkK0oc5euVP23m5nWgiaHW5U+UKLeimqbVxw5agcjW1ciVLMfzLycf9lp3A3E93KA0E+4434av
QOr2pPsVNtH3wz/4qMsEbnXosdnQlA2tqfnJBFDmNVN3VLmng7EqjBR6NSs8X5fT9A2l/9UK6RRf
V1D3GV8AInlmCfNEjlYXvMJHB9U0pNyXC8OKdLXW66VSjnuQkND6FQxB/LXGJ1MxOb0DzIZ7edRZ
w/WAd/dP7bbeze6qsaHd09E1TgG/ZLaPrzIx5WLqfvqhHCDDQOdRBRNheMX9hKbbyk0TqPoZVxEn
oAywY4ns0/6lFPZbsmpI269fqx6QxHsLy8oJOIF4kqKsCGMPBFfaWJglBOO8p7tXbtd7lCJ34fpu
1lMQkRTOirrQXMn/shbIwfWRQn0vzjX6JrteZv70lg2J/uy+FOdPQxwTNCVVWNU+CMs7Kk/JxbkK
8Tqyr1R433dd6ML1V/G6JJA0Mdexk8f3l2VRSYFZvzArRt+kivr6IRd9CkwC2/6RC/gI3fSPlyyQ
GsgViqaIE2yftH6vrJsPOOdND79i4CSO/Vi2+xT/IFZfJg6aQAqsLdFKpyYVBMmHPPmz9eqydnx3
1LTHetztXnaQ2WxX/HgRTAR/LhNwL19slZoZ8GQhPlq/uHyWnGO2ww8yY5C+zXnsfBOtF8bg2kQq
k1p13YME28MTT5u7ISXr285DaeLEzhzWRoF7t0YFAF+J1BtYF9CJk2gYfnmme0qcFW2IwvKVvFT/
Bc/BhI/S73rshLHQn/iO5ujEJf5fJi/qCj4G/FAT7PUC2fyZ0spJ/GUSFmJvpI6YWUTkXiPZ6agp
mMnv30RrQwOidf1A6Xfr7RwEIp/PFtPfj5OOqQEMbsIK0eg5IaXL5qeBLsm3HIOcXOQOKpkZzNZR
Dr/3IatsZcL0jbEpu0myn0ZD3dI4g+hQMpE8tqZDiFmpR0SWTaxghcHuh4PXt1SU1U1mQR/VUiOE
nrUM8Y7r8CjVAg+TRhcst5d/2zQI1aKhWEDQm8vVzyyWfgzVPHbJGjvmIr4yLsDvtJGWynpTw4Dt
LUJQDmJWPLxSrT35hf+gJBeX6ljpMH3ZOf6rvmOS7sSu/Kj7wSFFmEXa8ZZLoGgnChKk6/G0wZkd
psg8vVDbJijp67dzLD2nnwBCB+3Fbi++NqypSElolm9raihQsv+fcNuRTfIpKh1y1WXj6l60CC5N
KcMD4LYZRfU6XPhZGALZWmKB6E9OT5DciGByFrOLCXbjjQj0iiGqMNOoSbL7Pg6QfoH/IidKnnM0
yiZu8G/aFzSw3q9J0kIZKLd9K7heGmilBSRInLex2/uKUxIQ27hSeGiIi6Autj/NXQk4lnMXCiiR
kNxHV7kb30tgzsMOGZv0MIzd6QvBvkRniMnL4vVyk1VcrPkDJjffZROVTuy3hGqDHUrfA577cSOq
vZMc7NWSsxfCmpaVswmlwqgdM60BvjeBL7ye1V5K6xvCLn8NXz24ViqqlzPV/NUsGUHOvONxgr86
LDEzgNMn2HY8m48oQP41mUeqMxDHcC9hVkL9cKVsZf6sQijqnshxxACQJetToit6QJJAxJ+Rt0/U
6WuaSu7AzOLs0F2mV7fi8UgzeAsT3ou6iVIvKf478TFbi1/taLAYA2qcZCH8BMLHlkIyqsj6wS0W
TV4wspIUxOaK6izA2/TeCZawOBILKb7qRBkDnCIs+R+1EE3OxpZ7t2psSYxF4owzVmDOyTTgrn5r
WlMZlHJe1iwWITi5C75RV3LTBCoyTpLmOJ2PYu7Sxh6DOKXWci8STmcfLS54/Fjbn0vEUPzcMSLb
5YCG2K+CsO3Yz8qnXy8B20oNO1nN7Xd1idFsQ1WMLbrWhiRMd9khCIPzDb8WAX8KzbszUi4GrnKR
jzliAbQau62G8h/ga2E5pxTox1hCAwRrrYCCDs3RnDBujJpeGY8isXwVuY4js+S36x2JwK/z8wGf
Dnugumg5Yx3h+V6KnU5vGwbii5mZD+qRonAPn6IfrnSJAaXxyCXJ+0DTOpRokUNLAj937960tQ3/
WZhY+ZXbTnGeYfgFL+0xUnHKhLtPU4W+WIMP0UJVGBigsaafOxeomsTht3eP0ce+DRyl+vI375PD
0pAu3YEggBF6LmBHxEnx8p4etWVWZNJLfrJt4L4JJkGTteAecWo6Kx0/igCjurAL+u8fFRwy6yge
cP1FI0OkEogfnG65UphxHeYZIbnGpeeHmMhr0IZFGe+YuPVCZy6eOBnpB2ufP5alHVqzCiPhqNOq
9XiVhJlRVdyWuDeg+06Qb6QmNJAV3Io2q1UbmSW5g/zRB0WjbnpARQlZ1QQ1Co+MoPBI15kO1ijL
jjsOrzbMDOvw+dnjqDqMptly3ER0wExo0s0oLPuHR1Hb5z41Udv1ws2Tz5+5OsfX56WYEq0Jvm2U
6MEB8ZzxT1B4qmUkAQtaNPHDkVo8gcwS3wQEtR+1rUwOsRjkMC15UObam8bT6dFPQoNvKL4jMNQL
AStJyxsO6LaTPDqQo1UBkZu+O0psXTNEzpPIZJbx5zlV7I/88xI8W9psB79kWiMq1NPK8eqvaehM
6+k1CjhmnjlDw5VwotOnzllFZrmJ7JL1Nna6gQUdcDKeSyKy6e47spEO1nEyHL3CcFFoMRCnrJMr
0qTbTCRBoquGxLuCjxuw0voYsuGZ0sCLNvKmlt3/aCcgxUqzFyXiseoLuerMqBZo8pwWzpvbevVd
jYcgb370tOjlYbOUYnhQdz2JFMaCOQgbiyHCqLP0v0R1rlUcbv6zwwS0Ekgx4Yrmt1cL+rKZVY9L
wfxGx5BDDrxbisNuyeIptCJ31F9osCVru7J/0Lb3OtgU+7/C4oFD4ldy/7sC/A4Qrn7lSloeEuCH
NcGQia7ggWW+hfBvZcifl/F58hu4IlJzX+cjCOHQy+KIIEiaeYAFJfNkCHXCctFmdqezdb1RvHI/
WTw3NeX6mzRJv4TafvdK6Vgr4oWJ38ZLPkf/C1nBzX5ayytLRNdaR+BvkC+GOA1sshrXLYzRwk3W
P5upyVQqhAiomVAcyRmUUiyijCo92ufENncWix0zHQTxzuqlHVY0hV1w9f4E4byMSX5Kl/BCUxkB
615M0AElYzzV4VNWqHuSrTDKS7Mp7033tkrxR/aElrSWePcaK//q3wj3Cxp6xtipvx+Euvg2ZsnI
wIQFIYlZ3yO7pbwtVP4o5f1xHXlpej5qvB/Tdr73qCNebUouwJk3Ot2il+DLuDvsPWEr4tu/YFEv
PiBhUWidaxw4CHrxXNwgYUy+EIl3zNnm1DMxd7fzmpADfBACKp7GA6x3R4icQOlUhp/FoUh3MoUz
eDctrxP8j6qmnJ5QWGPgXCALRT+3SUaTgEbu3SQIkWYQ2fDpimKdpwff7TgZ+gGJ9Gl3dv+RM6GB
sHyKuE7d64u2pVvhOq6Bl+tUHXAJzm7Hwxbk1ZwxWrfjeA2k+J3l2Y/La9EOcgX1nOUXwdt5fo3t
LE3RSowoPbvh7PiRaJynRnD53SW70u0t1XU531mGW8N1Q0MW/Na8CWzLeWB09NTW/nEfgjiTqR8I
lqM9oifDm6bEfSQvMP+tEMYF8HTR/zdWJiS3zH37Q2YlTR3lLJdlaYg1nyJWKrkX8zvgqHSoMNrY
x7sK//rGjSz1PLH/zkQ2+chAMprc2J/hL+ZlVmTdSbSTPOYd8bRWSN10kvDAW2gnMLYc0+o5GpW0
rb5ufg4+mSvC7nd13NtKVS34PAsiQHL6Idf7UmNygn9BxJ8icvjeoRTBrKxPZoxReQDF2zug3hy9
Lrm6v7fwS9f3OvtPvZbYk4QAAK6JISJX3v7jL63R/ZUUtLwtcTA8UvcHDFU5LTZfEo40dcVXvjAy
8OTW34lhc0lLD6CSlcy2qxtQ/gysbCrhHB/IuTnVKogBfLc5uCerBe2YlxT+GJ5yD4Tsh+z/eYpq
E/ovImo67Efz2hGEPB2Vr+DQ6vP98JLk1ztHYzYMiL4gMKGRHp8Sxe69Ghtn5n771HqhbF3LoIBw
uaKwH6GW4W8Tmdyj6s1jioNB7NvwJ6rZZ58t6F4vKu9JnPUeGU2Zh8FzFpwXkA80ykt4FJRQ+LDv
qNy2iv9zeBjnipTWl33uFaoIsTOpRgbZjHmaI9tFCrWnaBtJcRpyg2T3S598iSEjh7oAgocyV4Dw
UYZS6BXTDhgRFEgpvZTpVQ1QnBB/vp1hZL5vFFDuLdpkyQd8uRpq7LCOG529NsaUFICaC7yf5qrR
YDt+6QPAhTwDM3ZmK+O39xtAuV+hlIbo5oRt4CDU7hZbEAN5aonLd6GYC4MyDpJ3SZOKA//wSCf+
F9gP8MyUhfKOVK1Dfz5gqIQ0lB/SCo9r2ESq45TyrITI4IA5QKmoWcU4iNy/+jZHNIuv/gU68R2P
YVlCjG3mXAtIZpsBwD+valkrkejKGRFlVJH2iAUXmzlZTBKKg9T4WWXHSh1aQgs+7d5eaRAPv+md
frtR3I25vXcCCN9uOh27RGLnm1+IFI0Daz+9YdWGBa8jcnMy+01PMGDo0JInPm61jqg+kglfWJ/V
6RZZ4ZWDUkGY1QKeMxlABolYaNkEJ4vtH8wKzZxuQb8MnYiGTgb8oqD2Kr6NAPC01PQ9iAdV4HyC
2XNxwWLv0TYSnzFCL9j9nOHPJaH7Sif+6MOqMBrN8iM8/QU5Wdig52qsXp3xR6VR5jxBRINWbnOg
ATycwELMqy7FX80lVzd1jQ3zuhqjmvpwWLpYUYQ45Pb0ImjNPXzn5dI++stCpfiLWP4VHoIrbmur
C7ecSCwsuFDhKMjDSOX0Z4vTDMIcEZqqRepMYfRgKXC7opWQpmb8Nkl+kM8UBrrN2lfNW7WKeDIA
eSaJhuR3+6h3L22KvHVvQfIfaNPCafPs+uNrLXKDMBb9srxzlwtINWa3PyErOJC6V7mMQiNKll2W
XiB0qQbLwyGRlGx5xfD8bpL0ohVtCKBrm7BpeDbqI8dmK4bZQKlhdN9Ouu/kx5gFO8dJEq7WLeHu
Jzz2AmAspCiNxyPY6tcUnmpM7wP1fHB7zw9Vs5meGSArLTxccmXQ1LTzzitBl2ie2mXn943godGy
AU6HNCzv7aFhWy/tkbyelYuClufl1jK9s7rm64BgwtX1UqI6rDLjjVhLTX+guxGtqJkZU4p2SPii
Qhgjq6qwyvpoXnKZ8bykMKApyo8KSaekSLgVmJXNZ9XtQ/nrGjRbWeCUxv8d7deAaEb+4hE7SUGl
mMpdSP53hgRyQZ0ZfwPi0BTddIi+Q1bwT6gZ7Qr3KsLi2jIxjPWjDfg6lIGeJOPzHS9ufJPLcHBq
Yx3OxImCRxC18g8V2sncXjNkWV63OXF0Nqwf4rWBFWsymkO9lhTi2BEirC+icDSttKu6sbU077S1
nIAaw0CXh4fyaLqNY1Nc5qcx+VHfmV4rDHupWNjQfXuvly4vNGUOXzoUfT/0Tq9m2dArOd6ANKmK
hwpCe+y8RFZDgCXvF3hVS9Y5Hwh0RaPDl0rvm/cHZtQeWRGZo0PcYje/jYqO+598qFCBaq6wALkB
GWEO9gYh2loLK06qxZR2tyaFrg5WhS2MaOoke5w+Tynl8WNBEYsn+zdaIZlEX/M7UuCNGnEYsMHV
eyna9pGDij6l3hLy+2E4ZCJZ4kU7x/GCtfs1hGjorpDQkWgHBETCkZdDrsWey/iZgqvqe5aXvV2+
r8+I1Sd3HlidWXz2PuATw3UtPSzkeiGEOCDUJtYaX70BrpAnVrsMEKX06MNxvtq44VQmfZd5lP1t
Izru4S8HzT30+GcKFhdPdmX1Kk5dJfFPGT6Vtx/S5FIgChdxQCsddmwx0uoJLMppcXg4V0JHCuSz
6vy3qFqvtipRr4UD/RfgDQWytos6HBWcelajCffVXfvgocqUliVeVox9X1pd05Faxl8u6dwVSVqA
gVyKYydaIN+2PgrGaKPrZZS/ormPTVD5TUs5/Pvnd7nssfrex9bfQHoxBKLhbgM9kKzRuy3j4pC9
XUEbPp/bqyPn5fS1H/OSb/yL7X+S1KnhNAZxX/kAVx9DHuNRu0o6/AjfKpmPeym6n2ykQSEY5hW6
EXbVFtakzHzXePpTtar9RabcZHv2QvvFfVm+wvdkXF/Eqc/rUOkzagoNHO2iBlhL+DT6dCS5kMxq
c9r08dq+khPxPClbjmvZaxHWaxqOIscnekzV3m/6BMqRA1Affj/frpobkawKQnHHfVoSh1NEbcWs
x2otRYfPmzqzT0aNMs5xEO902Bm7zVAXSVCeUQn2SgBCswb6zi0UpIJbSEA9UgGQ/Bm2lfwsEdzs
BIbu6qBNZ8POqa5vXjD6Fn79iTQLOFILh0McvrtYGwgGM3ROgyEAQrDdZzsyfeSvLQrk55tEU/xq
xWaLxmt+ZSb0YNv81DkpqGNgr1uh12HgoWZZ2J3JH3WPcWHyxO8N8O0KxBubiP4E1aRL8zqLVDfi
d09C5gkA/H8BobGRJ8LFF4G5OQoQjebo2DUycXuAnRRKgyQfzYhCKJwOGyAkx5H+4Z+1p1tzT7R1
2ENKwzYGjkZvFnHg5oczekTorLrxCChV3tNs4R7RVKP4LpgGK7YhXKJTh4T6xbArUopLTWtGYFYB
k7lWFmfQPBrlSocgRl9oh+svVahmqiUmwULwWh3CtUEh2XLutDA4N0czRMtGV8pMaudEdM2NyEuP
dKhbLrUKVSUo4yCWNCEgMg77HoTfRkxk7pAbnK2mYt02+YhOV6Jns8icVDCXKiPVGKOCQ9s9eC8R
IuMAO8wpUbYdBUkybnXXRBnf60Kj1U1cOi3GGSAfq36fGzSGjVuf7+DHhqhFave7M8UwVADN+PsQ
bwCoO5fM2MZ6ekVCRSToxnhGJPkSjGFMakRiNTs1FBI4sKy+xMRVQoUs3MEiYHXkhgwxrWDypjjH
QFVEZuzi2QhnAyls5RzIcqw+VglvRRuUy6Yr6zfjq4612RobF1klD/+OSBAsGU+NccBrBr7xuy0O
D+H9/3QZkToRVw1uWuQxw9/6Jj6NiHVA556zErY2wFInaXM3eYUdDT19AUf481U8Sb6LYkZiCn8q
vxET0BAsWz4KPYRfvRb84XDMQsXZB2YRQyk8FfiRyIN04zfXyc4d/8ph9oaZuVov9xlrbex+BpOo
qw7G2jdIZS1LjfKAgJQJlDpqjq9W1riYtAVxWIOfAm/PBZzGRIR5plQwCfEo+PW1h7PjY8NvE268
WxvSC2ZZD4b2qLdarNT3dOfoEM5DxEG6zZMA5rBPFl6AdxJ++/KFBiWJDfW1xRL2xtLgkH5Ssr/x
+mDRT2K2dy89ppOAuKYTzQJjgpns3Q95A7/TDLqj/kxKs64vRp31pULNWyly0RZw8HqGgwWFfFVo
8hZYPkAdgRofDG1d0EZODc0obV+KuISJbM67+vlTiDM/iZ2LIQhko5JzqmF6fKBA4VeKxkV1vm/q
sHtsam7MlWwNlvtLhv3wX8JAUDjYkGPhG70sixDIfpj/V3kr6ZiJkySs0OJhJKaOOdod9mH/uVT8
WIQgxaJ5nExmFh7fphMwqVmXQNJ26+HiDdFexqhlZjvDOcKlnEaiM1tbcQxCOkfzlFzeDNq1yzf0
4vSIgnLm2AgWZwyy/eR5BinBv3vwWhmoNHW3FCAv9NSvu6V6GGWEp3qM4rjiHLIXOGtts8mfO4fe
uv3oK01OHdAS+OGhTEBHnekpQ5/IEzYhH62phxGQ2y/yw+R+sNEOSW2ViH92ieLy7QezYwe7UwR9
YINNUmDapBOEXiyz5x3EnhdpKmCtm69CSXXra4WPMN7jBYQo0y2PYBBDPR17Hj9BZQv00A16+i0W
2x6T9EpsVZwJ4wmOdgI7cwASdq8vktS4W7ZH6b/4KuI/Mc6I6HMnxAr2Okuoo0UsfT8MBJfUOpCk
3flA6PeRSRCOAqVe+bDqKRcACaDFp+JoL38bMwuGvUnJdenb1jqK8iCXiGcP7iMbOdgl7KVTKGuk
77eUB/Otc/IMaxuPrZMway7w2cMr6ZZ2zHTJ7Jns8Cpj2nWbC0+yMJDpAbGeW1cqETISoWRu5uEb
u38+vjJsAzVnCrCwxafkTyeBHW14I6AL5oZs1fsDIT8w+TVTpVeGbE3Vd+dRmzX1MGRaVk45MILZ
cIIsksVRQeUGIWFl98lSTImvtoDdiXcy8v+o7rhTwKm5xJ/BDFFIEeAHjAOqIEyfkcpof6oncGQX
IksFYmtTEoMasi8P0rpuWaz3VB4ifYG/lmHodObeOyOCQVMNGpSVp0P/qXuAefkNSQzpHv3I+lX1
r0XNBCazYX7Z6jMYFW4tupJ0aX42mXTEViJw/5T9QRFA/qEHpAAyDSocgPeFZ3/qPLieJcCIvp+i
gjDCJNBCopvEMnOQz5ZPJYiciUfzrajV8kqOHMT/+EWReXa8UlVu2zw3qSEB2ONUEzIvUli8V1uy
/iTbU8TpEoJOHyLJ++LbNNU5e1GF1GBam2cWQrAZE1Be8tecS/aEakIf4D9DuEy3aFYXfbriUzJs
9yGOvcUonYiUwED17rEc+wVfBhntjO/SH8SwdsVNOvRr/fjiACK58r6og2KFSE9bFE4GnIkU4THl
N6XCLXITIiL/UvxkaiDx64gWi04w/DBphjD76Ml/A8fKyEG4p0wa/+zlQRLQTd1KTGsLgeDGJXZ+
UP6VKebci5WdmAjji4o15ZSKvuLOINHJRK2hFowzVpP6JfVBscy5oih3FQxOE9MV0FBWyQBD+sTR
5ssdCw1BYOd3P3PyUoqmxy0Yty1Qfz7SWDTZhZ+8S56ZkhjYtb10XZKhb4K67/MeAmQgpP2HrqhH
ltHW8l9AF58tZfWjjo8bLGw1BwwLeOxHa6BC4CHXkTgYrbsYXgpmvkL46902GFVgopK2OMV3dXtl
/N0c6XS6xh22/JUjiOC6SLCM7MB3MFzmAhBlRhFQ4JmGdd2mYMrViukcAnKKRBAVmV8KUOPIYTgs
NkVhwTauSgkQ+eTz6g/yFgguwJiLUTP3RF4AJPfXyy8J9wX7y+E0N5ivayDg7ot176Sz8LdUghOY
+tkvJcKJOCJXNrJ20dwf5gbwVLCv5mRFpgMMS1NWdmBQckxs5UEEE8uoJ203L2BRWa1PWPPHqScu
axOF3YLdI4HBxeD3psK5J6tinRvQ/B07WxxRK3Eng9q6lLQwVHPA7BVz11x6aXSQhhTqjMhSpxNI
eagvWl1EL8nhJpKsULhuygRvlAbU/obonSNSfjjtfFqOUpjVBUCTNqHk6YliqINnaDhKcoCnpTll
SBauGz7TUx+RY0XCcJScT7xSCORQ2dshZW/YepTNovUZmnH7q1bty9w75u7Hd6QpuOMkh8y1CFe1
Bq6HHQXLiEe/KI5ssbzMRVDaOYMUcaKBEWtW/4vOoguABb0JIokRnOpRfkLk1532MV8KmypeLgox
1QMZta2K79lHrpcGsiXF5g2+FVz1XNbUpZ04VF9KARnbam9BGfNa+XepVm39wzJNnU0TnidmZeTQ
yfQs6D1EG4W2/ISzXcT+OgnAnAubFNrqoTDy3iyrAWX7sImor/tRo/cAcJuyyL1Ts2vpsuCQjP+d
NnPO2ZmcowvFCu+N8vfBwM3QSp3v5ICaecST1CQBbi+BfzfsTB+s1gWzihyPfb9A9u4z2DRLqUjg
ayNRDShmr/4Bwe1+HGaMp6vhoQbYFpL7uT4kFWrH7BY61gqKtRdoumo+kj/KtTgm40Ls3u48FC5o
G4MY8mdzyfsZwnfkBABXsnn3fEyWMsZRBlfhrAHWCVRuUu1PMp4K1FEbgT+GA0KVsIhBJ5QRLj5q
bhF9a7L7cyMnW7Xy41fnbz20VJoOXK3XEvUXfcweHGei+LYyIUU8ZJGFU6LMZzM05kvQOMDluYb/
WgydlMdZ/S9axWBWRmFK2KmkfMdPx74iA8V4IWVuiRajRDmzHBeaj/ydOeDKQ0wKBn3dTvHGUYE5
nHLOzZ28lvOksBT5Sm8RNe0wtM8K6EU+1XWAX4iWKEz3Fpa3a/hEXY6ctghotJcfmGiaIOVSCZqF
SNP5+1HI9O59la1+IKujDmsRplyifObvlYwplfBJp1bEYwrXxR7Zf3BaN/8nelaOA/DNevnzz2th
uZo9Gr8wK35bOHrwgmNzJuLiftyEmaIjonejr09F56is3evVWIwiukqBV2XQa/3keS9Zk+CSJ6/C
yNmEevtL9rxrz+I1SyqgJZrFDMX1uHlD6/4WKpe59zzqnwsgRbWpC64WRvAKGjtFOOCPPXXHDKWC
+SIbu3Qe2806GJ7wOkVBJbrIhVa25z/jNfkjbzlxRey3fUQMRzoPEbcqNNBwJFgCMQ2zJTWmHs2l
etfDeYibVnDYgXktI5+/t0kDY0Sg0yzf3mkgqgXiF8vii4HRvy4UJdgmQLsVRBfW0Wi3kOrCgtTc
iF/fQvb/KuIyHjS8nd9m+g8oZpeys7l3vH7k4e1bpEucU3JUp9MwMRpiM4fldd9/9vtpn22MdMXE
gzIxRNIeqF3iaUMcqnmylvGjE8Dt5JvLPdyqgC4U3gyD4rY1g04Y/7PPmLNhYFP/oooE8nngm+NO
XKf5ygiS3+QZkrXISQ3TLncg7LA6BeGi5TPgQW000Mg2xUkJtDrDkpNFIodUdDuzuH6JJeR9qV20
t0EjVBWZdQ5/zwqbZVON78nd/+du8JvgmdY5i7UkITwCII2CXE1mKlWn5aEx5XooGHjl1z3hIltY
xAGRx6jYHM1ADxVnlyByN98VA2CVQALdeZSjO9tnHhJ0d8GMCIOz/nezPoTycqo/aOblH45nrQ4O
Oq1aGCU1v+yecqjIKuqQxmQbfhDpKT04VLnhnvsBwEZ326z6toIuBt5UHSxDn5vNonlm+Yf6B4/o
TocJoCWfZm0f+xzs4duHN9k+9okZEQ/a2nIyzDaGDHi94avViXoBKKoV6et6IppQPtHCE4R4A3v5
1oEdyn2oZLOo9l+OELDB7tKkkDRfy4FiBwU+49jtzH+wx9MuRXqV8vBymToBZSVigh0sWi3ir6sH
Dvf0bcUzD+ccU3iDip5cFbYUBfY/Gkf/JBXe8GdaVoAsje28hLmCYdaE6LfHlBSJQs6XvNR5rdtL
4twVUKbDa4cPIAyVpcXepDCnaarKKJUxjkvVUchqwkinI7ZPfNiFTL0u3hLNJoEH47okSgzmm5QS
nFpN1yDzvMGHE8Le2ODDEXBhVdBeZ+1zv969B/FRLt7pKACbk1J4MpRenfKFVJ47JTPaLt1kcTjR
zTmIUqOg25vQJEdrjCvF67RLT4eij8SE2UuxF4s6XwNoy2YxJRZMIgGZPsQ1+hO4BKnz5wFLA3ra
d3F7ZIvJANlKbvWlWBj7WR+g1NydMy4+vM2PZe+28rKtnRN2Pr/9/1cDRvDqnMI9HSOA7wsx2LR9
yzdf+bxFCXnvkVkR3ASwnhk/lqWsWN+42uLO9fmbmfbmy4+yAhrkyIjSxYzxnBcdU4ZXew4d9agR
nLTwcGgn+L6W+2v+NWkUNcBQf4LSAEuxAD/HoQG0xqOtKPi6+YLYUTWP2HDh2iyqvDOFSr9nbM1O
zk9dBb3BprLWzy7bquPEbjcXJo55WBJozza2RK9xJkXkTd9U8v36rUbtpMKf31aoIPAZt9RC4LmZ
Wc+Etd0WCksJQLijTgiC4H5ijOq+ibidPlB6urw7l6zAq20F+ZKc4n1AyYrahjnx/UM0SJduUz4A
EkBGjV10d8mERvkXlaBeaGhNghE9a/sa3O9GJ/hcy0KMM92BOlyYog3gbenBlxtliqLYYFJF0KLE
StKpxCxi7kyHqsH8qlzFdI3HaJ+TWlGGpSN++TDdYhW5PkZYmfmgDnH4ad667eyEVQgEe3WuD707
tArH1hD6o/A871xMsCJnX2WigDzGXhdxUqsnxbNrK+tmF9QFfZDj6xYWeNh1Gvv+BvoVfW7bPcIs
wfgVVedw+b5XMjfR6gYIU6hZ09+QaMgYNPZ8XcYEXWkNtXVwKJR9M5SlwKmVJ5Wb9GFG++vhaNqq
U4tnXkXA/WSXHrduBmrCuCdIvhrg2sWFljyWEX7qQR4j9GEAH+0+hGj8v9aFVwD7+5IQJbnN8t/J
tYuWDAQ+WLuqhGEX8aJxcUC0Ngxdli7KIlfp/KkmjI74pQly8unXreaMmzH9Hsst9ZThjEsAmJfp
WQMWDUnmz5EM6Rqg9TKmnmJ8QId+rdOx2aVkxym9WeigjhEb6l5O3RKskA6PLOQ4li3+hRMPXKVI
vfcOwVwwas9v34f8yV+amxG95gjkoxkWms5nvOCLONGV6otlZQdihitO8mNWYyGxvaj1s9raP03Y
w4soqd1YteVGS4j6iFxxkEv0s128eg0MlfyB8LlZfm/44hUz/MGjWZDgqQH7OgtF0Tzg/Mqwr3Lk
W6MkaRjZFle3POGS2eUJzZlcecdEOIUDrmvr/POvdqKjGcKyoWK9YaoxrGlpwRo3fKQWZ95Qz08M
BnmI4LDkBBeIvldJG2pIQSBlh15gZtPrvroUePNPKg+/7e3MjXSma82Hr73tbg57H+rjzNLi//T0
TNHz5o+n5TxBPbQrwQRXe0v+io7Qijkls2NTlFtgVcB+z1CcG065SoVJRkuV9+UCRGNh2Me3F7C2
Jnp1mkpsWRoR9qyW+ZVACpGDwEqKGyikxPvbGZvyjiduL3zHplxWOJQ5p8D4HRC2gwRPa5utwZF2
lNlhpfCc2z4Kys99yFbWQWd7CjM19fNIYchDOUxas6tEd1BbH/0fyrEp0Njtj4z3ABlptBEMAVgu
3zgJA6OasCwff3D3LbwOsTqWCqh6l1EzwpGhanAR/M9P7kZAoQNxrsL/Mb4DF4hj/9Tmm32Q2Xt5
csSMaiDTbrA4ZJ8q1uXd8SvTirSaD3EP58lRkb1WWQMlUnhIqmtI7/nSQJpDpEG5b2ttmVRuvtTo
L3gngmGL29fvm4VAyTQmi1EC1KMtWA8POA/b5zWSPOeWE520LoXI9oH/jMp3RaFYcjKB1MtweyLT
bYrfQ2VuABlj+ZYEJ8opx8FmPOJ+D5Z7nF+RatfQBjlLcKHgikD7mjL2b5PBzIBEhwHSzWNPUTAY
v9zDtDbtN9mLyRZiA9xyUaCL9PzWgIshDzAtFKr9IJ3rNb652w7jLCjV9aL9X1mOBCi5h7lx2jIz
A1N6BI/PwV/Ncv72dUQOkKDLKnfpfDv5hurdatAWLHnkwekfDOdE/wxwAF4Dc0EKXLmWQoduuFuj
8B8kerff0mG2KRSAjp/UEYp8Icvi/UJMvTCjZ9/d6AV/TfD7KTW3+LdziXNkX0G3NrR6OkJBXzqM
Z05GoNDVZ2IC/sUmUj5oq2v4Vjl/2Z3A9aOJs1rOa59D/X9iLBLg3bl++HdXCAkrRjY7H2rCR2zJ
EJ1kdrBnUVAjQJdCNC1V2x8YENBCoabI0MrC8UyOesHGsdr+uG2tFIm61MOUi7ZEYhllFaEGP8Qx
PhXEK0t6C3IhC5Vib8XYi7xVXbGFazWiLOJLSu38hlZzAfBsJNJ1WwWBgkcHItz1RoJ9Qto4XaPe
RlE7Y5tGotjMGQeED99R8jxRMIIOEi6hzlwsyYxTowtxUlzjS2vL8WrerwLZhIRTkVPp8DyUKmNl
QHBaGxtdl7Ojp+NlQasegjrCNp7b7tMXjBXZ1HkSDE0JE+zepEOLVG/VgUTOTl/6R55UWKYg4oyX
Ug+hLYRtKKu96AcIb/WU9LMapJ6M64vDwDZ3kKCveb+ImU6arULD+nNiLxmQzkTEujdPrPrv2jln
wTyu4Ea7OAyns7uwGHz86Fc+IupH0K3KQ1ofJW1v6u1XcNmRCcDYgVNM4Be2Oc7hEeISPKbMk0el
7EaDEYL8xlunkMublJXhog0rQRcEFcLWic8y22XsSwMV5fX2rN2E9XgsT73QY4YHeH4/jHcBJe2P
tDwHXl5v1/cME+y1L+xE3f7F8n0kUbwYO/hZ3aWXKjlcvaZpo22RqBJvfG03hT3cSXLq+mhmKNmf
wO+YIZ3S9rIIjQiVw5bSvkdtwo//FHOOZWmbwJnkmbquE16BNA7Iw9ezLVmF6rCQEYwSH7k5A76Z
x+9QxVh7LB9AcBpQ/Kofv/LZ7JDSRt45YljpSIhDN+6wIdMIhWCxzroxwI5y7Z7bNXI8WXwRC3/H
BLFGDWCUnhSn9S9V+eT87ognqHF0VwuunHRTVQZFlAYwccW74fIwkEOlMlTZYKdp1GeSOJ9zpZKb
tW7GTNYkl1D6D5sWYegrfW+xFKPUEZDGaCzTUJjPr8VUInNR5+afQ+kaeBLrbk9XV5K8JzAbxtJ7
CHHh5TWq8CfDoXM3DXlVSfsid4gJEXnGziGSlasYVAETg6i3OOC4nM77Crppq+YR8c4D/cfbN5Sj
gezEIy73cCc9S4qbYwm/4xes0iGRtfPgka7kfnom1tRl9WDcl9ixOb9MbSBhgZR4UdJwyDS+gR7d
z6Eob83vqH6b73r/iZnIvAEZVm2BcMTSb4RC6WkmTOzHgOlcC2I6nn1iHZvT1vmJFcSL7OCOLbAv
WriXm0WKQTktE8mCefWJqstNtnsMaOTAR4XZydl5m/314Zp4gzva2/NJkWGeVRBldv5fwJZthzi7
vigQXYMr00+oYMqZWpCm4f1KJwHh8hPSM3zYHH0FV3cvLFZlc/iuBS2PXr49ZohHg+rUSuuPynWv
APDdGSmhy0uXiEMlsGCry15BZR+WPvGHGivfEUeqf4ABoPpsFT4rwPEy5+MnAm5KMwsdXrNyTg9h
em4E8ToBCS+lwfLoVfOaOlQ2TuQKwMk8zXmY+hA1kXl/BKT4EEzQ9CuAmQedargWRz1U5zj7LYKP
+M7KNVqsejYdgZUT+H3f1rJkqwo6j7i1XbWqDOMgClw9DRUyzZ2iiF3QcNQfRsfWBzmz8u2PNdHe
Iy9dy2TqD/peQGA1wMdysNale+eG5+CkQgOlDY6aWhiaSq3Jtsib/wKAabC0hiCLSBlWyOxMD1aJ
ODJwqYxZ1mAlVGdurQV9Hu7iYfJ/FaPH5jhqLipPS2G+6s/e+hbE6NGF3li2gJTi2389Q49mrc7M
zy3q+GVOQ2D+I2tLfzHsb68n3WBnCNv2GjS+E5Qe9+HS8wRJBqNTznEKeJGSY1W443dawLRAN3ph
equy5CtV/oOAjQYrectD90rKUdDVTPkqjH/ZKJKpCXlYHygv+z/5hNn+zw9jLMRvJOZlae0A4Y5O
wCJ94cMQnhUDAfTGsb2+H1/el/ct/Vrt/xTCcl3k0s88m9tIMv/v1RynusqNJs6jpV1haL3NkoG/
IciPUCygI4GBQ+fobUe9kaY5MZ93q+hhPX9me/Olm7E5y9hAFnBUcVyM9yE0kSoo7wlzKx3JpJvj
dGEYIf+TElsStn+uaceBFY0sn/4jAAdR82H6rN55z/XG6QT2z4cxcyNaPtLHOnC1/hs8StuO/acD
X+v21J2RnLLR3rUR6mQJH8sPuMQzacrUjPJTZ65I+7oo65qsZOC2iSYtk4VGFWFxymTxOatFnNxC
y6m7+azmh0MJDOkWzU619oQ7EOo5e4q/uAbgBWuNGzYGq+VTne/S4Ec+3atOegaitlPvXmIMfZHD
UFIJprQeGd/fdfBtKcmSDOqgXU/wT+BqpexAdIgZqrxEZO2WZptqE0tmg9y/p5d8+Mdj4I2QoKit
MzJBVeDfnRc61Ty4JZqN81l5YmYTyJgMz2EhVvPUXmMhWFxRCJ7gpaMFsoO6F5EiytOSeVVIEXCO
F33hXjVSHquoK+D5TzLDBD1QVcaPetGU4qjcuq9Iua+1HEawZZfX2GiwI8n1rlfV+0owHtngoEkV
ivIt2QQYY/4PtZpEAqAHq20ysk8NwUkP0myWI+Z8bIzODf9pLDbDQqPxQbWqTrcjLGHEyQPlXj6O
0NqzJBoEbImBOxHTCCiXrAz6tgI4sHtDju5ZHNmpUy+Jy4lnZiT213xBVmb4SUY+kqwzqnyl2hhj
xkVJK1GjBCW/UdagK9zxjGmZC5uP++vqMW2MrWOcA+2pyc4QZvYN1llnZIezmIWh+OpGWgq+j3jZ
42MQNRYG85vfGIjKwijb1yq/Mra9/RBC079L4L2Y7KeZg6jfLWgmvfoy/tdtKtAr7pgpkav9Gvj1
4sEFt1hZIrb4m+ZALHxxh5kEJw6OZp8Y8/fByvlvjUd6g/Elra/8+OpeO0jHmvzlvMYis9p7Lq0v
966LuIKH7Mkm273VnDWT1jqPPhDKU8FP2ZiQy2kN/Qg6t0v7mipljjBL2Ygc6IDH8hd8YmM7JcTc
ARS3zlUe2NoDglHBEJF/5DvCatB+rUeVScHt26YpqrEvz49q7JAHUSG/hUnQVUDF/A1/Dddr6+Xk
HOI/VrUyNX6yhBg8FFZ7te7gmUQzzYZ8gKNP5ned0vmlzELILi+lLe6xSxrYJ8XieSMRytp18JdA
J0LvVJHyhMvBZfXef+XhFpPKWevNIUVFu3UtApiQK7zGD77kolcbCc5nCh15k9CICNrtwaonUipD
ZNa1Qi5EQAEW/V76XRKRz4HRbzHjoNdWbxHbCZh8Wf1VjkpY19LKOCeeXWHpi32l7KiS3b6K5vkX
Wv0BFkqlyPJUcOP8iT9qfizQ/n3kYAC08Pj+uShQev8hVjLQF80l5Nif6HvzxwRzwlCT7CZycfH6
zpUgUmCU1/cEXEOI3i1EhC3+qxCURihlhsuW8hghQlRjSPA4f3IfNUj45nrI/G5qG8C+CKqcgtDW
Nj2Ub/EViSuUkoWyx+Q5tWM2U4LVqFz40fhj4+CCUgj9U2mgsGNBuD6cK74gs6YwJnPW3LClt6dY
pwn3mgCCIhR9AxZiUvc7Q3YWHcXNedtyo5wOWOjmkKPlVYwDY2QfdqovstznRUoj50RaK84VjHBk
0S+nWC5EkJWRynjbPhJPJ4WlgPtGNU9LvIz0zR/c27to+esEPMgCAo8VobPnR1vaGCyU9EUzG03Z
TElx5crTwWQSdmQ7aqCG8AOrFGDLrMbdstjRuahTiZAs6nsiXvzUc2ZrRCnXES8P/s+r83wWxrnB
oxujRGgprl8XlnOPjWB9UA2gJWks6gm8sU8R8LF6YOYS7MJONb8lT40Ys4y1NmnRGmKf7L0UcN88
9veAsrYGr1DK4ArryqwozUDhFYxNx5kET2yYFJ2gTKCy3p5jFMvJM3wD+N2F8lgrAgfAqT174khZ
VHtjAaXcLkqQ9l9G30MoUwBFLXMx1NOsu6Jfw4VuhiHrMe1dpqaFlTK7ZCY4nvQig6Au8JGpY3LZ
6ihq+u1ar34v4cOLc0dlhioSoc3bNzFueLM1ZTTd2G2sWSfCBa6rI3Q3wJ/7vwC4IJjPQDCV8i50
ZFvuYOSD8m/9ggWk9zjACBT2YQgL2qG2lCAql0W86yU0sHzilh3JRpCRdRSt+BOubNff/EGuAFE6
y6cNbIonwO3sb+auwqZGBbvfCBcDK+49inxeTWlIy3+2vttsHGL+XydRm9oQml6HDJcP8bVEqMQa
7Pkof3Ts7mraBhJ4Us03WYn2Zv6UZYiSW5KSWQI/4VV8sj1kTrzKFRzNlCnDYsJsyRfVdNNnZVmJ
5Oo8XEpH9lcnCaFADs5aUPuJdRDeTNF5y8gagpYsb5+6lh0ocCB1c70r2iiWKLA+5dQgX2hBVZN5
kT2UHGScB4wT8C8O2Wbk95B/hFlcBmutRRPGT1FhTCoPr88qDO3sLVIxBVCmLWJG/PetIPuKXu/d
Y/1M6WzJSSFphh7Ir2m613FhJT17ErKx5gqSwg85rbel/kuaDisJsV9UaH6tE5oMCB2c9dGB3Xek
0exnnclLWYsEQ8ey1y74u9V59AYfG+8FYMvQWOFiTVEuKpSQNaLBIF5eK93K35TExG1JNQ/5fx+H
dHPl5rsaapuEaq1JCYqT4BHkaTh4GVCIHfkgFpyfn0rqZPZnoFt+XDhyLaJ3Hc8cUbLA8clmfVh3
82y8sRV3UeQKnypJbCmBNQLOXVlzKGEKiWF7FWFAHcK/dilQQv3Y93wKUO2oPyPyWktsjVkkG9Th
1YrcUktMKmc0PE4jaUekjlLo5GgOdNeq8YvMFF6X9Fpgsq9PW3RnINoEdqXXFGKs/SxYQ8jSRTbM
z7ah5qAMjxofDjfMPElbbQZzaRlERkYi+CMG/XjG0ZRNM84f9gLFNrPmC5E1UmZJ8B7Unq1uXZ5G
ce6iw4rrQIs6Q+7XtTJjzLANlsroBwjkmFjLR/QLf6odshh5uGvsd3tLF0ofEUMpAmML4YB2P8jP
o0Ff1DV8aWCYKIe0+h/UY11GXm7+O0lP8+QGWoX0ms2g7RM1ZEVKYUKjrHh/DK10uOX7V5mpuBGy
yE+5qiWtnH8CotQeleNXkMginwHKnbTeKoH3sTdrhFWUnaMIVSelo4eu8rUHQR/GL0Ri9CJsHBvN
ZepabeyPhOaj7NOCpy7cP9evjY84OxBabex5eySrR8yGkRAisFBh2xcPcz8C9XT7/pxeWNg1k7Wx
W5DC6KuInRFdpJRjJ4eHYxNwDxNFfJNydcBb9A0sveIiOYMpahgsrVti5lPJiY9p+a/9IULAJzR7
Qeqvyj1goJgFWoNncurv4+S/ApkdjhAQEpez/lQaCzLDOGU3qV8XiYLoLtcaHaMXsUYCqC325i0R
9j8VkpOTGBzwF6XAKW+vswqoKXq1KvyS6AAn4hIWk/4u2AyCGT5+GGKW1J1+PVSoPvFJZl0L6yNX
omlX2WYWENaG26isxJbQFfSvMYWXIpgZHAmY4u11idxfQiJ0lyA+m9Y3ag2dvIXRqe7IUYGW+D+5
LvF0MsIvkxVQuVeYbqYe7Jf8KWxxUNJQ8SAEIIVL+2MWk0mkgefgHEprz6XeQkxLvqgbJx5lymLF
FNLUSjD8+8Nyl6sEjjtvE2UkVg71WhfynM2uEKBbL16+19nJa0c9K46UR9r3FojOytR1XOvqlALH
MHi9g3Jt3rY4G5z2Njai2J0zYWDnkmgdgIzdIoCsH2MWJ6PPhBScxUK00BQBL57Mw7M1hT987NDa
B+KGVuI4Apufmbb+YULLkirls8JMFsiK4xaSRl+c6q99F8thpb+xuCSIJVN9mjM2gbiefj5R79zl
cJsStD0ZY9qdoxVpzimkr6KjGkaQLiNPcp09Mlh50rGdHvEoYhi9vXKnzbQg3ZU9qcy7EUbhKUqw
Zbjo68CkcnZf5ihXIJCQpVmm4Jjew+/WNT2NyjRiFUId1uvFtcom6MUd9y5NQRduzoutjqOB5b7b
gw2q48Ba/34ssf9ehWs2Ng9QktyI/6sRiVs0s8uETchNc3fh18EKOVw8t3DJ/NXg/YNvcA/RI/A5
tw5o46Isn+Ni5xw0oAupkiYi/DTy6linfScsiS1QlYk9WdKe0JRKZTU4urGsJszkyfFoq/aXo0xQ
WtprXUDDw82cv6HbcHnKk7GC+SD57DmxXDU6TAg5TGryl3ungqjVistnlgUBN3SaqN1+7DDoT60H
mK0rs4Dm/PfmsZX43NXONq6LaZNPp/jULXyrystFWutyAPF9shu8DZBmBeWHx22wGN5rlhzk/RCh
ZH2KSnVDNWX/7hQ/ZziV01+rBa3tbagVM8EtI/6b9M/DBlSh7RKFNJRL0eTNM25G811Pa3BfhDF7
C+o/p2ACI79mAVz5DrUl9ZC0Dpd4hw1ITc8N2XM5GY9+KMLOOoyN+wUTtCv2vL9VpE/TYHdBZm0O
Fi5nI36kydjIBjTv58UKulNxtMwaCMd8QvUsi1wRLht8ZNFjcq5F3yvy8oh4cQohmGDi0qIBWESy
1ypYf/kHVhQziUPyJxMCrZ9JP63pBbnK/jsPSjIKbpmmptLP4G+tveSOvLrqbyUiBpL0nArz1vzU
lM9WJWN5QRty6dXMtSXsm5Jr3XVCyqdwLv6JDkfGaGSNv4L74ef6EBLtLozyafOhbMSAa/CmVlaS
uah7/btqfsPL6blFTrWnydCoGzXBP7ycoL8Lf3FZkp4kHkGE/jns5tAEf45HnDqVCv5bVl7pMM71
ZLpTLNyYFgXZoO9m8F/S7c6gZ/118+0vfMLKri0HKyqsqHBe36PANpOQIxU0YTnJPmF2bVqHCZhw
V5ticY6z41YKv7JlcV2qURJhB8D+o/vObXc8Hzs7Oa/9LxtUQvo83WHfZDD13f3nJmIV2DSfcZwm
0HGyfJ33q6ZymPllgio3W6Edn9LsKS9CjA7m0ABP/WPcuL6Q82p4IWSL3omaTm5cYK3tRxnte/aA
7QtasCb3LLqJPIHZ3v7S1CQC/zYj2IEQMSp+WDKUgsSAAAHsTXdWI3KRKlzn3Ih5d1PSkILGIeHC
G2Q11uLiwyltnmmjtst1kuoMnIw3i9CI61lo6/NgUXbxVZ/BBl5/oZaIzyC07mo9XnCE/xKvRhq+
tg6epIOEv/NlkU5Q/bU8QhX9gsGtTV9UQX+n+e7HjHsQm8v2dfN8Y3kkNxe0+jllf4ziReDq+7mE
ZKjDK0y7XGKdC60OvpX5RBaWwkyTL5qMQB1EvkfPPKdmNfxf8vU12qaAwJWN7hXniGXsBlGqBMPi
+MPi76xRyZhGqO2n/brDMEfW1A1/eD0YuTSbCyr9rLyCFpkXYY+eQK37ZLlmotgVy5MFBBEAbBsM
4ryzboXJnpU/5BFQHuVFM0I90YQu4M3Inmrl0KwgPImHQQi9dMdFoDWrqKdyjlP98apj93KYZraN
EQPlNHNJncc5+rzanfkP3gX0bUY3hx6QdLzlzLwXWE0zLO9CyCEmts5JMXIssdh6h3APFbdPJLbu
BcEEOZL+LZXZCEwFqJT9UMy3v4zv9MjSarUViBwAq+VR8vXgLyytp9vovmPKgpC1Z2dPuT1KDKIK
QZ8rmNS++AsSA4ImUVajEvYmAThujxm4Cy+0opRyPiNo1wDkDLernm7EoOcZc99tUrfJg/KMj1iU
zDAWonDJNrGoSqA5u2EnunqMHdBfU81X57PiYKNZi5RCdZrogvsXg9HiuV3hXkNXD/we10PX9XmW
NpMN1PPf6fqnOgxJCS3RaIHtGwF6vpVEqZzzX2wVcySLioHijI8gfWNHmBb2sMciwTOc/liN6A56
1i8VuQ5diKW2pIzjELqUNu7pPK6AROPwfrtc+8+peL3GQHHTjUqyh/lTr0AGepIZam1XHdKWGkne
vptucH8+YvSiRQY1x/EFemhNmCXLQbR4QJK+ZmyWvTDmzEAJrHLLkJdlJR877uDyUnor7snELc1r
FRqVAGBEnFNyOno1e4as+rT6MfAi2rLmSV1XHCRAnIs6uBaeYtdg3sDx2K0tcJSr6GIJ8EKj84lG
+CBmVHo1DJEd/uxmpna6eutFKliX+V/FvFLj9cdV8zClgH5cFgR8uSOxg4bhxl/XM6HxOnNyafyK
BINW98LIMSmJLDcfF3YWuBDOIviaex/N7UwAIdgwzg+xn2S0jmJlBLeCNO/Ui6K0ZGAUABxq4R8I
xE25bLpvmnE5AazTNoHyDqlxa36y4QdpcEU2IPcyhJC+ahJALkNMzQIw8dtLRtxzWlBdzDyYRS0l
T9LKhmLqLn8NHCKw76wsRFoCXOJnqtUEwhqcisA9bSh3R8ax8lvLuw4woHGlKTJqIf6nGj0dTXf/
9wWAzClZidj9vtLxR01ojLCXZKSE0V7Vplve/89F0xpz8XiJ7Mm1Niik2QZg4Np7yTMhgfA5ATJf
LoTtw8DNAJVWm4Y+oY0qmwoHui2Lph0aOSMVUj7D5C9IbuZA4QuUc3uTwOVxadE3SBhwc+9a9UkT
a171YVzYtYiR6SpsZkIeHB0wBmDmBFomkGD6/jknojKCFgmoYVowrH2nSUUgX/1zgnjg0MDRGI9M
HvhhKcp07+7+k7hbUcBd0J+1+TjHDKmGcHDiMNwjK1nAKJbjizsz316+qduzLExZlAis3fE6sDwq
yP08hq5ZD9ec5IjiDA0uRML+pWllOgr+87K111MPBvo/7jahU00y0MlkG8+B0fc+opRvTfAyafPF
T1Z7R6e6oYfYyubpw52/OsqFuUl3+bfeuPoRe+CF2ofHrRSYA25R/Z/Lgyd9VvkE48eXgVfSn44Z
GbkDIU+ttV3cvpptqv6AgxW4/AyXbblUQTS9Hc9PXjGoMa+UdB6YUDdOUvdLOo6y3N8BY4BiODNt
eLcWB3qxDkHW66/nWEmOi6wCOgPwr7bIEcrQW8NpWlQbrdSo3gIMdQvClrijS68a0p/QMhsmD5BG
MnbRRL5NTEehAFxytmEU6kR7TT3oZ3SRZo+9D1AYCuGbN/pQWx5Bp5teLKn7r9Q+RfJ7uYu4ZKY4
+T0LnbFvmkbgbe/d/W1ImKXZQ1pXDEdz9TTNE/zIGsv0jB9Rjg0N6OMpInaSHxL0oIDZp6Jq4rzT
Ezm5kDc0ybJVauCLXQwOJl8oYZpZzIqKSU5dTDtcjsbBGybiPKR4yAi1EH6LJcqL2O8aoZ/CGlY6
6ca/OuDgFG8MH689vFjD8hmJ3jG3kHdnNwjp9Kpa78gU55Rp0mQ3fQ/hxpb6iVJbfEIXxxospBfe
heGV3euDeskHOPkWsplKmcwsDXrSIQTvx6inFdGZcX6yLr1UOom5q+zf4Ebl18NLtDiEn4ISBb0O
u/T7YdPk1f+RjAMzsKHVy7hGbU+0R8jSB+z0kiGvQsBJaCprfAm6166GyOOSMPuSV21dtjgnWNu7
nBNl4+kken4k0ODsXnvHyiiWzEdqW6PWVdB3A+bewnLIzTdAONteyvwl/Xl69ZyeBaCVg79Y+gS2
BzEz5aDJS8SKxqkEWjdEbubsbKkaIIcNwXgmVnt2C5Lv3eklOeUKUof30dFrvv7cA6tYZdCt7LGW
lIk5Zaa2y/vLDqwX+lTZaKoebtN/aVc1PYejozKFVag6/snP+xaJe8GZirU6JjpWQiNRZmB4xV3l
ANDK+d3eal0heNG0iwx/uA7aqNklKSB9ae51VS3EF5RlPkewnG7N1kLprHvjlw/V5T7kKU4wy3cF
xrir2ClwRIju4XMoZMjl+znQvl4qMAeCXTbaymZiE/sNRKkR8t/NGENRvmyiFkpLhuOBhIDVL74V
M0CNNgznsDdiSR1Wz01U9LWuqdNLasKYvxQGNwf48R+d0iNR7qEkAKHkWywhV6qHiim7gLF06XFP
h7OfZyjZTnfvvaWQNKX9qzpigh/vY9vIZxpH0Kbz3q6/Smu/s5lAU+pSc5ZMXfSDg2O2C4UkACQg
nR0N6E8d24LPCBbKZ3vQuFDo29T0D9VIM0JPSwLWKtsDJqjdrfYcXZqUEgRKcHE9Z2QzR5cyGnWV
tzLkHveg2HWl/yTAV6cgCq3HVfmQF0gyI+sMoDzTMP/G+FsKUr1FC2y5hlnf++dHA2mjajQ9d0DJ
eMqF04VFU/4JxbdFkfzDAwhhBW6x/Kdzqo1+5qgNVRIP9uS8zxEDZdFr3wiPv5eI3wqC89gXwlNf
bjEWfNeL1zPecqq9tOr3bcto9AW3f8HI895gPG3DKV6mVBIxtjZJA7OHvt2x3KuvWvU3BkU0NTyX
s+Ifg+T5hNEKOzvqiQ/rbPIhk1KUqGlr3wHR7rSB1pgtdAR/s4racG6WAEH2TRv0Gkl2M8109tGj
AziVxtrl+2qnXgnmS/N6jXkSnHrpU6OWoU1iasxR2OKw2Q2SbZg+CQ2lGtv5wEwEuEcZ/qrib1V3
tMUjrDFUc50mhoh1Pr/vxImwP6gEBJx+WyW7RMu73+Oz5He87TWLJj7GHCaDMVFIFhae2zzUTGkN
ToiLkSFRZuZ5FcpxpxyC1LMF+h94XS9or9DS3EREtAyp4DqEMLvjuzWbL/1T1PmfJV/iEs+t9pcU
ayUO5tVvo383wM2zqZXBm3MUItCyRK5SmgUGxzcMukxIAD4Ve+K4VhpGr+DCFS3vy4SkbpvrsgUz
+nzAd2jA2wtuf+Euy4rR47DDEbtgiqH33dtPvRKk5lI7pdaJKRwCfPsBMIgB/OwhFLHVkuYYlGPX
kf876TPsq0vmfoMQ9TkIBo/nJsludnI383tFRBsQN1pTBfuHq+s3nNrs6HpYqpwB1rxeMkVY1mq/
hAdPErHH/peJbb0wZYREk0Rh7OKKPTISWqKlSFwO7H2htypbiGePrbaBvkz2yDrQPohVNUMbw99L
IOW6E4wcPEPkqn8J+APg68knZDbnhn0uK2S/WYYJLOAEDOMJoTxLIzDVx+UoGFIDTrb7+od+qfJM
zc7/CbCh8LLShbW6mdGS3wnbCuiP7TNz6uEIx7dxjACn5Vyj6+suAhxP0bJzsdzZ8a+0YyitR+Ck
DoHsHw6KNw9We+fBL+wLJi0zRlNVWi5GyZ0X+fWPCyhpWnAEnR8JPLstqSbb7si6v+Uqx/WZjGQB
omYxd7vgvlekCR2g033iqae17oSNkPsFfq9Nm8FDQw4yD53pVkCIt+5jetJ2dnx5OnEaOTDCLWmz
1JJwDQxQ98r01oVfVXsCdljat55XJnHRe7OUd5s1bdpmU4XcR/8vLY0nvaBZGytNj5gUrnTczSQc
pNjApiayX4yAMXQGGrrxt6EHZqeUC7XPMFRIOw8uLYxTWV/WAfQkOu0eHurLa5EP3Rd+Q5o18yk3
zAy1SJ+HElh9qriNWrhLQ3qOsQ9dM02TbBeBwvBQK9GKHvqKDCz4eEzaDE+sfoYQ90UGqItPDHrD
FODphk7V9co1s6WVSwpT7wAedPtMjC8E7/v4oacKfcs1sq0gTwl4A/eM3vVyg05I4Z453Fk/ur/r
b5hm0gZU2NClGFmQFOL96Pw5JRFYGI/GjS2Vuv5t4CjaXnY+5s1uYaFEHLmTWdtdOkexa3EU89U/
HLluduBTvpbh/L2xYjWX69yxuygNG2u6so/ktPaKEkW5BCF2VMRXqCGvQmBzyucyoVlwB33SxT8l
w2xnW5b2oXa6vUfMQy+0noDBuXtH69Xx52J2AUI1u+WMPp+T9DllXb0KpBQbuu1nQmU9A/o6prYq
KOEEmhiZqwxa28S+uS2ZuNdvNSoIk+QYcyNLtRW7X0ew8n0YVnzQOeq8cXXdTDYOWVDXEHRQ/5ca
F8lAjdUHp4XcmrJIM7XooeR9vzSZfR7l6L4I3RGf0KruYFVTREPWuvH+hIAY0laubNpMMhAFABCh
pGIXYSgqUTAvqmP5AFUDD/T8A06J/HhvGiLSpt93G1cK1mbZ+SGkbJI9b9c0n0m3ZoIUAvwqv9ih
xJPQIHXvJ3bdCgT17TytKdhYEX9cfJVOLbjumbOSzIsaYyp6lZ3SvnMtQ7gdba8XeVxUew9sIJi/
JDroPN+EAsdcS+vls8IagzDVWmx+amkszzlPActfyDmV1UBu+fCPiRNboGWZBmfnLFfb0PaBl7Ra
bC+f2aPzkx4cBpODzcU1XVo6U74qLtVmxRe8c1O136wY+FxU5yHYIkfMwHwrG3BXAj2op87kHO3q
FDEQ8hPkXAZsx1b35PRDGMab4Oxi807wOEMCzI58awMRY8yB3iTmC39/qH3RxggXgGz6xPnxwa5O
DglPLz1sWy2wCaipWjrz2A9JDMu95ZJpV/P7yJTKl96r4tEG2TMv0ykffxvhj6RxjSFQRS2MS9m5
/JpcRfIqazLc11rlf4KzZ4GORfrwxxydIx2QlvDz2t5DyzUtFBq1+R9iJOjxzRqbNw21xp/BJsPn
gbiOQ8N2ugEEZx1Q73eaUz317PRPLFYWbDosgDY2baVQ+XuQw4UxYCrJBmAyEayn0U1kC+GFAzn0
bby6h7AGMahueVj+cchskh3mW2MKs13I4lS2kWMIO3XBBJedv6oDDYOtt7gBU/e1SBIdWC7eq+og
3e1962s/9yDSKy79TIWGX5B/VxpgMzE4uRM2Dcd2FMmHnpOIcYx8hwFyGcwQPlCHwOFdpPQxfwq9
JdbxJEc3nc6jwMBQq/wnb1uHK2Q3N/G6jRn34ZWfpieNXdomH6SIKym56D6KoWkcB3bltZM8d9D1
16Ne84dkCTP8Sar+wtptIik3CwPd5rqOepxUG9+FWgRCrR1y5gnPG8CQ2oyfOjdipxTGwdP+3LxS
/3AcRr/XQmUKe8spbX8jP7kv1iJMBmvY8FH8Kh6ma6xPeEA+uZ6atscycrIMGbWGh72cGeBZcRTC
ruLmVZwBb2EHlqK8jaFXyzELDFn3dwOHiyaWccLN8lVP9Xk8Zyuw7PY8v1XZ/7e0JmuUaHLMF9GY
KmcavBe2OtH0iGINqOot0iXzK/lys9/MSKbiTWwqtY21u+f/zyu5NU0kX7eQVDsvLnh9OQjWxPmL
Z5aD0fpEIooVJ3uPparwPixwxdxhouWyEMBdGCxE5E/hjtq7ZQTQEcEjtl46Phc5JOnUJqjbViFk
NYJVYSCj4uvelYIwZjtdp5uE8oJI9xGt0PDB8uFyhZd3vCL8fYWBHj7HRDt4n0GP8A+7Uca5wRW1
oovSEDvon5JnSfUVGRYAZsP9wq1JtXW7kC/Ilp/JYsGMI65WtljO68n2PW57DgJrECwlyDBHN9TT
/4tggkmjsXPAxibL9W1yoyQpXS0GDZ23Yfmax3V2o5N+VxYG+kGM/XhbUPg0NRsH3yrBGyYlAXuc
S1Tz/UOJRt57h4oHqmaWi+EEpp+VGgEC1KwggZl0NyQMoaymb5MqHsAP3XMpT41z/AQn41WsCfdu
996gg4VsglP861WB5XuMQTvG14XwRibgTZ+Vp3ipLenqSlXzvPw5F5GqMYzQV3Poh3lXoFE8G118
wIUfaOK6glqyE2xE36IDcPRtRb9aqYAmFmx9lXWdXyEGUKi+fH3vaShRBPO4hZBLIP0kwOaLV3+2
s6ULQCR+wvGCTsFwRJLvl3j3kwKgpYCTQ7Opff8RP7pbN3KA2ksJu70RQ9vLrl05+4M9b2vcDOC+
RxtxmdFS4hUkqdEZ8dNmBe0kC5sjQDWpaRRCjb4iuMb83KnmUI7xfqb5KucmZ3zIcR5f+7vr7g2x
rz6bGRxBXUzjwxDDfK1DT9YBaeAvbU8rgcAEWw7wnDLiE8PtCXbcmg+Z3yWBC3jgoktV0E69WPTb
YLRCHvPat8mAdENooKKmZmXYL7BfUlhbATPvdvqqd5j/rQ5IwsX3hL4aA8NVRnWyNLPddPLeSjg+
wbS4HUFDZYT9qhK4MFm26aSQyppUAGgkg5jiCL6RCQ+koGMU6nSYXZdbOBFLw6MKPa8qb0nKx/jB
ttoq3yGYTDynVsi0kVxQqcVDD83CM3NiichlIzg7fI7XyK5R65l+DOptYL2gP+Rd3RO/cwdHp2yw
Rd6dhPleBjjZtQ2SWBtpuExLu4pHWk+i5AJthaRuaQiXT04C8CyyG9sZmdTQxX1740WJnHVTtbHG
fDZVhQEy2NrBi28z0LnFQP8knstHwnD5RoxRYu6QpqBM/m+erQf8w8J0Ct09SY2fRvQLUWlp+s/Z
FGzKTRiqasRAeRxLKBtDRY2KmC+7mI5qgkixtYsr7OA0USfS3X2Kl1ZHdYW2PBVvb26Uwak9qeis
sLX2BMPqip0/oh8garRxSCe49SnCOZBsmGAYxgo+sCISBksJU5CJw1BH6lTO7XEsepN0bsFHeTXJ
L/wKlWI0qxvG/Eb3TthIcmGBOmMKaVc4C+fTCe75aVJ1+okid/i5MzizmQVyl6Ezv/bFLQHAhIBp
zwWKqCyFNhj0z0SrjrmlENq6nNw0jmUDN7TeUbEAyq+mdkfG6RHAp4R0n8kms2eFYL0iqTkXgkhi
A3rnoaHmvGKsw6AboVSmnOrBf7muI7kV4YDgTRvaZg8xX0tyqiIWZiPT9aMm0dxdUogJA8ieuODW
gYp+Rh9rLvBDMx8HAvENN12PtPd+EFeSzdrsyE6vG9gHGZijN9beG2xZ/OEMtGZ78OvZS+tmIuqi
astdOEArb4sk5yCe0XgbwYiSazEVaF522ojP1aN01yMzxYcQawqIK/M9TQ6O932N3LynnLhv+Cmy
egC1GuoaufmatAriNjNEoG6aOn5zq3TJCwppW6uAnA2RKYITHez5pjx536oakxJkTE8Z6sg6y42x
vP/eaLgqxTu6pQG6sc1i8ZOq4DzGcP5l2BNRde2giLt7ncS84NKFDvMvElYginepOgiReO8bgktu
kA3CvvVBeB4XU7pMCyBcgb9phifNsw5tTUu5WzlIle2zRXa/Fngir0Z+djh7xAmFTmYRXJbIifX1
7Af/fHtlKqaCa1OpbMNpG62SGdt0NUnb/mLpyJjSm0zHfIP4qfpzh1W/5harq6WlQzkbnBuA/fk9
13CbxFtgM3MyYthGzl7wPt+pxc6S4UwYKVGJtm2XOHS1ZGQCgW3Lt/knucQrTevUAFqiKUx7t/M5
OIokErTusgHfLbKcj3J8Jy5/c/v2c0YrhfiNtRu+JCed4CJRnKgNsPfqnGgpPbSwbqMC1LcyoYUB
jJQ9SN5SQIzCbYF7a5NQiVCqR8HecynaA29RO71OTxLbxtmRnjfRNLBKo5/eTADNwWQLIXxPiJgH
B2I9YOf78b2YFTTqIQ1slEyh99HFrblQ9QNLCkZdUAzoxqS/XlQ3t7Roc2kW0KvGxCUdVwawa2UE
WvGLecl1wJj/iTFjlzd5lqX7Bj+Tf0PV1MmosPC3i6hniaEB9rFkHcWqMl1gjvjG1qs2kBbEzBVW
Xm5OXanIZJhp7lmjhkubbazp81PV5UBRFq190ml/m2yy0v9hEcT/5FJ4Li4etY0Y7Yh39OGId46t
C6gi2+9+gNojjNGzfIA5dZiUWoUkVFwd9yWE0MDFBb8mTh69c3LKb3Ezg4Cw+j5fQE5Q5t/DmqFS
Sra+MAPv9XKjN5mz9jIrp2CZ13/tVrwh01yoZ/ZYbBy7JFv1fY9pe2nUFP3sOmipppVXKt9CxVD7
SFgaJYVGmxBbkey7BAL7Jd0296gonw+Jpey/0QEDYn6oOidUJBtSMXy3qYcD6GmqivO8W96gBEZz
j8Nslu2JcX8lFiK3IIAMIMhhdy1dlpG9or7VMhv/mHKa+JZxi5V3hxtpVCiRLwjreOFyKBugUEVv
GaTULl/RmrHRYCXSJSHVn4qECXpGl042Z2D5IRB11+fTPVVkhIUvRQn8YoNRM1gUQCTA3iW5dIQ6
e1ms48FohMFjjPVFc7OutKmHV9NpUwUSYvaQAw+varIFFPJzkrhwCTkv3IRxOEakE5GrbqbAImPr
MkbuHKa3kP1Fd/XFPFOLBshpeuzyiaO2k0rnmadTa8U52GBHgjINYkHMB5d/x4v7vpjUh5erQ+AT
pKMWMEJ6/qLVmbcN9bXnKte+DJuc6yR1vqtGNV4eEP2MHvV334NxpcOtzgv2Fk7yT8dk/Sk6UHjG
Btw55fFGuXcpMHUjuxs4iC4LFtfL1hHzY400Mt2iHDdggQcRqMlnvBmAp4PyMoWeosM7F0m2FjQq
KMbc5EnseYf8x4PPt043+iGG0mqmoJQSmWGSzV0YlyyrykGUV4z/y6tYHufksCiW8XCFmPgfL/0p
JM9q3LwXO6FtpRlZW8Ez2xwuqrC3BWonp+KEE2euoUqBA7ithLsexquwn6ug042x+96MHb4ndAto
A84QFuNh3T+KblwPdCW9FjQqgER7gAgi/Nbpr5pBZM0tqhwTR2m93mxRaGqcvco97Ike2LwCm6x6
1J+L2MXCJVnuib1yYhkXGKEg5zRmqir0ZaJTdQTMKONRb15XZG8Hfkwf5hrCliI1m9tUkCSS2b9H
rHBqNnxMAvFOXHGy9Z1vERch3ncV+rLkUDjWrDjFgZxi82OWtYSq+GGQSQx95fLcxTjxWLnUlM4Y
0h9J/KEXX/PZuOn8AroPhJqXlw0+dl1QVm5ztKkWLh30YtHqQ5C0BR4dj+HKftov2nEZ3Slhz4Vz
m2wx+X8Fy/5XesYj4mzHze59GD7JMWzTLI8r0fBWN1gYHyOGhL0+i7lJyTjnviTW4/ElpMHmk+94
Gy/x1VqCVc14RbnqmPnC310/ZwSaJELEeyGu6hpl0MRqtuU98kBvssLNahGMALG3G3BrD5s0BAub
o+nJ4uG2ZjNdchZDZDrGsyTHlBrqlNBwF2OLMJR5DICTCGrU3nkd6u9kn8QuAkXYi7Z9NdsHua2n
ewGug+WmA21mO4Gb+Q+O5fx6yL3Xci23GOpI0kdDfCZ4xhfU2kskcbeM+QgffE23eOuI2RlZjJIK
ddlzwMBthi72xvnVqXuhgSQLxmWPMjB//NUijxXEQqbNetQqQjxRY0aRmoHKCqQREueLZFhvEqud
Ze/yg6q5kFd7zRz3+jMFZstPNJ1G2vwB65VvoP7pxqZpU7xxgna3Rj3hLkxAfum4tqekwuVAOMIv
IELvvh0FdnBOOoBmrgnv5e64GEeUZWsArLnRCjeheavBHzbMEvWXHo01rGE+mJ2kxkqJSTj2jUQC
HCWWr5g2LJbF9pMDAWTRxlp+ZZCAtQP3MmX/DL1u4S+AQscrVVw5mU9VJUy2LQEBed8wTFcKOiSU
D4W4GnAQxuAGbR7K4vSUke4pxsdyjLrwTV+1RCWEaFMkPYol3XGGASQblgjYNUTJWGOHhAIyBmbi
QTUmoB21uYbJHV8VZj2HC4YpQxeD87U0L0tyv+P+tVoRLf3FBZO8r+CQMeJ6So9xi2aloIuVh479
Ir2wQ4zYL8WvYhh4rya+mXk8yagON/YSoDjb25172dO1tbZaZVXa5fH3WMc5sUhfawi5B/U47TZ7
SHc/rprA9UHRt8SrpKxd1YWUY8gmQRF4wFvRo4obj6t7GPllFCbEsoBxvPCJtD61yNcHrWgloFVf
zNZyNoliFIomwJD70dKyGG64DRy9qErf3bxIVbOvBkxVB+lhXTy12Uelp6su+KP0thol9dASrqGX
Nmf2cR2c7kvCQ8x62Y/N6OuHa2Zo4agecU0Zo0wNy3ZfOfZwCcbTqm53bsmFfQ4f+ES9/PsAGRxg
TIEVTvz2WmgQ9rd7sd68xUkDHQRpNcpv+CV/f8hX464BIPMWanQDJQodluJouegPU3/F+NU3bNY5
v9BTzUJcX7a+Duzmb5XVvAElMZVzfJinuk9EFUr4LPlDJn45TuaQbiTSxVyiwk+zmVke/fC2FN88
vS4iuMeqiVioT8OWhvdx1g3tjHf24sdKmc7/271vgi8PmFR3v9m7dUV8OTqwFN2fTL7CYlNAU52y
vVHqKQpvqXxZMYXbi5IY8IhMrVHIabmpFI4uU7P7gINXleA87oUjyys46kuczxO9CjQs/vlzJvnN
19m03m9ukc60nv3eBW+h6iTph12v4B188OA37qIs+k6EnsO1NaLnVKkoEM0Ay+Iyds40o+HxqYvY
Dj81VYIEUUMJYPAB1702LUylhOr1QDOqT6HX5LTkySb+CoUX4EH3X1NPmy1AFj44kGIzWA2RDpRq
gkDZ6UL+x9qwEMPV9cYauoS9Sr5Rr3w5x8YpWDddtkSkTZASyb1yUeO9wSwDAkcsp0Ih98lfGOAK
0Pc9K8YrIYMmNjXZLQ/EZYYBNi3sHKR9vwFPMjV/TQicZdi6FhUrDI/klqbwekObQsN6OfBU6q1A
/GIU4QQ+eFytuXIt56URe9u+yG0M5SBBOfUD05wndlOE7Giai/u2zS4EzFsbIr3Smw68vwjQX7Q0
vnU5NAgnnbpzvR083CPz5bZxLisMfXgbdxLGphggTfZbA+nO6rNf+HoA4Ez1H5vIx1r+NT0fp5NT
wLW1QuEaO6j4N8KeVfrydWnkZQC/Kk35U3r3Co4RTLMAn0blDtuXd0PxhPIUBAIdgh8adnW75cXk
hIZgzYn2wtAzi2HMQzS/WdtpbWPe09pmgS6JWVGV2jXVv/lwdQYuiYXAVOLw4DLFI0pyJ1xLrqss
WGWIGz9AgZ56vuaruuv6+UBBSH/ZagcKJNv5wQC/8mIOhTR9gP36BcHfBg49XbMxtUTp0ZHPvqXs
5TPBBxSXRHf+7CDf5HnNaHzHtmLoS2a2gw2/lT+SAQmMo5hJse97IMoD0VAYCLX3gqMFT6zfzsCv
zfWXk5df96JReq/0U4ls75YoK4+sw0exf4GFElwY8hH+EkY9PESww8SrAhsGwQTZdi2vf/X9xEYa
ON9IJfVyDKJfTZY8den5TbhBS2BhJpuVlRrlskQpxn9FdGCNrC3tzoBvXkv+Hrvy5PtnwJ3jZBhH
i7qUZtnLllqyPB96HSmiypfQJZoN4EWp0/kdyd5B30rddEId/oLIrJqvqXLs7pbogvYxDyc/aLMJ
NnICAZ549of1eZHHyjcaOkPOsC0rDBPk1BVxbtykcdF8HyV8voix34fG0VZBVvD7QcOTu7bOjJwf
h86baI2WeEbBkkWx4NwM79PbViDut3N1jHqe4zabVOWSjNCEYRgYyEx4dTGQi4mdpJGRjAgKqeFd
MKmu60349nca+YZ+Zn/PwJC2GZ27RlCCbVBVs9CIfNFrQmZVKhVMC+mR3TAWODr/I2XrwXtSrv8B
fw9RXQ0Y1nUp9FkQU06tfsZogEnK9Wh5XL94UqZdoZXfRY5gs0RAeIQGR9xXTe2RiWbRwYpiolwI
A42dtXtaH2FmE2YslJy2UPGNqBJcOvKC+uQ7k8/FrTE4+J6iaUqWosvK67E6paulaIhcoZeGJbDm
sKiQCIssCQ9jA8bSlawl8A9rwZ6SUMRFrZSmNL6FjvRWQZgk7L5NpPIB8yBpfPwf4TlH0852hdp6
Ht5HKbI/VSW008XsPqTidnWqrdTWSl3eGSN2LPQ8HLgmjsXt9dSF/87M/d/KlZDzQmnDtjtNsqo/
yQ0FuDR9GnAmNQtZhpq3EeRgil4weqPaCEWUE2/ADUcqKArYaXkjcX5jrU9CJM57kIYwMuDlNNOZ
J3mw3ZRnFQAdu7dgZb++gbaTCQLozWmeuUb7DAosNeo8rpTpXrbhhUMKsT5IGD3rmcJARJb4rbr5
fsVqeXobt4z1NLWUBA0jbE/0zuDsrB0XnUhLg/ijHxYIM826dTI7HKymBUGTOCSxY7ezb/hoEPuv
18MLlTcWRa59m/9skORhUGp4TXJ0LBhOWZeExQMtdincQmn6eQiM3h4KneuWDcZjF7xfLsWnEL3u
XgjeeCzCYcTobW9RRwuA49JYM6WLc/GoD0iThoQqRgpn1j/xBrRsnvnQb4OscfQSoGovs/L8Nttr
XAoHkTbZpGNBcBrYgmtp4pQ0PITQoW6wsrfsOhn3YVKSkuUE72T+QHv7ui5zIrfISM9CbxdV193h
d105zlT4meGEtgx9K1xSxzCVeFPrEh9F6zWIYW+htdFqqULsngXHXVzkXNt3QvukNwFIhgWCafKk
OTORsPftbh82wGXN+KzRQ0SgEuGqvI8kiaBkgbwzc8hzJr8+ZH20sLZB2GEnzEpfGyKNGjz878Y0
sbnEMfW2HYfgzRBLQFP2UTNCIVkoH/MrbY35kqznchFrmSV0CV6XS2q505PmZf/I3FQyVpNfFT31
NzMqD6/vckDD63B2JtzWv0sHOCmOxSvsZvFT9PJ1izpGjspjCvH1DnAIjaM0kefbEONN0Z9amjwj
LX2vfBkI8IttfpDM1xuK3LtiDRiUVrKa9o7SV9AFVXuhFCm8FwqCpBcC8xQ681b2NMDJtvzrrCHD
L++amc/PDCT5+36eE0CbTi8P2aY/sJkJ9XguilImWrOV8eSHu38eS0n3cV4P8+MFRP0r7EiOEGAY
XzySNm609kx9/fmAxKbCyAZMgBCY44PQy78vYXj31wBFBL+lNePFie6vbTmXHJe2xzlwrOyd5N20
whCBNviSdfjKbEE2W0jGQspETMYEZfIxobZeeKuQ9uVKraq2pBi2q6TJDoqKQrtHYcQPyQ2RHJ8g
1hV4yGDcwNhOG6k7rh2Z8sZyfzEYQwwsUvbczmbfLxfJEi1eEQZKNWf1DIWnWzoDD+6Tw3FgqyVM
0B7jFa+BvoBJc0nVtfX23/Fe+92CucVYhBTgixFzCmDWCd4SSLpjPpBTVqDoUBFNi2B4sz34Is3E
R7w8RcX774uevQfC47TPoNkB0wIBxdsnHBYPP1Nddx5duh3vRTDw2of5XJ3MSlhFiDKiHx40JY12
XhfWpf+ALs7eopps5dN1C7NjI4sqaNWwuWcfPDjSO4UbOH7j180an4z/YE7mrOXiiqxvgOYJRrXX
wFxy83eonGbws1H79hRP/D3AyRp3bXRv64DK67/w7Srml47zA9TYwctn0Z8tePgJrpB+WB32h+/N
9G1DYfNw7roio8BFSnubC2w4F3ZtTmYXFyf6ZfeHuUacs8Q7THJZ2EC9aG7jzsLw9qvKxsVM47rc
ob5//hF7NfGbqRhBleJQ06fwg90f5pyaMKa53ZIvSuTv+OVy7GrjhZ6Ow8QNbTrsh3vJtJhf1K72
4XQFgaMjh8w8xN5xFLk9BbygeZF2xR7LLSPIurTqK9Qgt5EgJ+mMQChRXRyr3t6CFGiSiK/9KIJD
hWpmACI5E6AyR+gvRJuEPoJ8qhVj+AO79Eu0sP+sv5XcXtW9oW52MhWr53nbT4MXavJYFIpDIyej
zzuD5HSKVhcPTvnGr+k/KMpni4xLF/IaI3T2rMWCo3ZzuUKDv93cvYGIat0YkyQaX0Eh7dgD9kSW
XL/xXN2GVPyU/AFW/MeuAG3wRppbvU2DtdUYih6pbbcocfHxDpjlikAVJu/gYYuYdhZUDkebGqxB
tV9C1jUN7j+dtEjf1wHrS/zyCWbKX/rHXYEDS/JJaUS5QR9Au2iZ2lZMJ8xaELsBGzerjiM8YTbg
JvpOxqKJMnPzzsVPJTxOcxrgpKeLfeJaytnwot5+NgFK8l9VgruTWRXJOSsXchrFCe7a8aoBSQdi
wraW+/3VLg0VhjdZsJ9FhMlLkX/yinJsw80+ky6feCQywkAiaN5BhSDXpTyLQfvpUe57u6QsAmkF
d5JFP+eUEEUpxBySZbvChCD850bfVPpY4IH0hcBRU8+iuypaMDZKTCF3EtMPbJugQ2ZxvWmIXy2j
jdpcZm0Ftrj8pffa57NfKMPIt9kcL0kj9VwALdnKhiEPozXiYcu2NEWZRBXQUcVZc37JcS+g2FXY
qTVxJB1eYSG6ypgzWObL9jmFG8ebjDwVF4cykpWXrQTneW1MD4Q6JCHrmhoOC2M1vhZwGWtUH6ne
yBxE2mlOax/0LBFzq9+SMoKqqH+JPHJyogtQCQSLgQEtHr/jGF4P08yziTId2nQx7Z2TBJEiuQUJ
yogG9A3n0WDCdH047iMMwDd2NtSp1KeUVF/vxa7OVMXNZ9RhaMac7YJfqFop19yxJC/kVD67//8v
hcOiTH/veA9+CnPVWyPmS4gjN9WMyw+yJECBxJnnTuTPfZlCT0UyHNw9vhJVY6q+3+d/61Wv1kut
w7r7Rzi8yMfKwIiyIRWJTjyfVhk3m2B3mr2F3IguvUYZ8zCENbYeKebI6elNrRwnN321mnVWa+s/
KH4KADUhdD1+QF/YUqV2nuUAEcqvqAbwuOBiy5pYJ6bmcOvGagNXST4PjgbpjmEXhvkJOfzIDhAn
h1NhINGxxbGha8C3IQq8LSsRgFWrM3GlYmByIwezz//w136AlLGI1/11SzmeON5P7p+C6WfzIMCy
gL0uP3iKPGKpxpoIHGgZkFQw0hn2KgsS9PwZCUW15jjjaVFtzGqmDLaBUirlN/78s/WaJOssjGsT
wk74NSj3fIdSSbwKnJNF3cGCbC94Eoul+/Lxd+sN/yzPwEYlXrua3yUkBw/OU2NrFvrOkqB7kh8f
qo1AN0J0YsS/0OheaiLu96S5uUD6dFvihZyM0MRYSRsps53hWycRVoCJ9wXAcMhnKXXhgxvYlNTX
/fflMx4Mi9LIQV1F0aftub38VAi+Bnfv1xzu/W64F7AG0zZnmAHEmlig8hJ/aLRgbiZFtpFKalQY
k4o0HnL91PhB5t4ebvPytbbeo2F+gJRF+5Y92HgG5tK6QQqY6MyJbwxPufp38g9MvLZsniAJE06F
oPkqAHOgaLOBkYaf/vNuKkf1RTcDtyfkjwQEeyfgI52EKGjguSZ9V7ySYalXFlC8tkS/hZX8Peaz
JvbrKpxH5BSix3Al0PD0bo5sQ37gvfvyQojlzx0S64V2zihXcReBIr3qFVZLf5SRwD0RSolpS9JB
yWzhiz/3JnKdMfxpt3zClsxZC0e3wU44Xb+2RAFZGF9ljsi8bBDRX2gX+B6+0AZZgvSakfeCzW+E
uAianmwbkuX48i3u4Pr00k9cKC/SYfHbWIq6aB/fErsgVMiyaYa1K0Hy2Q/hcf1hhLZnjOeOAw8R
nDdyhbdQiVB4AQwvUzTN5oScWJfjhVuDIuQr7ZNSOjoonSPcvjp7Cpy6jY6wLYqHO1tsi1dRVa7r
/7ejIlpohkZAWt5Al48tpS9Lv0fqW4NWWfuNtVsVMQ7ebSDZb0e+FqV82+fhlGF1VWTfB/0z3896
rHOa9EeKNSvlQxksGxKsXPs814xwTfecv+d3Oks2/mCan9WE0N8RPaMM6SsNx+gFd/rhGNV6HEH4
im2jlBnvPKq3IwvTHegnfeczaXwJ4qkAVS26qhDG4JiFkBhw020XI4AuZeXRa5g3r3vukoLQ1et4
MsrZs/jCaU3+RclQ/WUQJ/2joqOA17RDGIu903O5OwPuYbvlYHNzyhw0Q0yzCj4z0eAxNL6gnV/k
v+HN4hXHik5PDDPxBfQWaaG9eLHXkmGkclIpHEo3f/kUI3xqNZCU864H/2/g1K1aVP53WDMXAKP4
DwXlCVRVZt9ltmkg8Sy5Hgj+11jM90CztglEOaFqsaRu7F9uNLcUUi3naausVuEZ6/2pHzHPwXic
dexqWPbH/NMi2oAtCn/T7Rmt1ukr08rjhtaXAkKziLclfGcGy7lATlyZqvyTcf/MGrLOSlbEWwL5
EKUus0cNrsVh6w+5OMq+TAeCbqKUm3RXd6L9hPPAVBn3ftt6zhgngbjmjmFVYLJw/QEaRu2RMjP0
doea44fr12loxvSwOCBRsMcP/aDWBAlKTtwlaLNY9A0WpekZJ6nIff2yDWKGSJHhKQBU1+uWIoiF
7p+CveGYa3OvwV3AmdOLbCP/nvHlLvNeIOChZBGBr8kDzqTn9eaya8a2b3+mgH6e5t9NDefAMyBt
XUZiMSSh2In5Ev66+mbXF1mXzl6vGh/CVEo9kEPnLvNoYs8LgV1ROcvf37cU6VoBVvuL6b8csZhe
DyAiG7pWGBPT8b6NJn2DziK6O6WnsemgX4iulSquHCVj/WGbn8eqw+4hBif7TGA/uwT5T2d/msvU
DygLJ9uxjY9n/r6a5p9Gkb7qksD0N5zlDWBeB8pgrlYvx01BE5+JEtTXGV1+3sMfwG9129Xd+B4B
RxU4ZQUt8bcDYQeTDiifaz3Q8ls6uhFpXHFdov4vPqqiS4mSJ52A13bktBQI1NVkUYmNSBKJZnYr
t9OsYXM2cSmtCr2T7EFy2RbcJUOXMuHNkTxbrADAsLz5UvaCqS+j8jmG7cLYN1p3VIdeqEMtlVGb
0B513u8+7UbtjEzq6kfuo7kO8quyoAQSgIPwSXJJlVSPsTHyrvYQSUTN+rbwS5A3QvjbvIrFvELQ
m3qjA+ZvX8QCxORIBbRvT0PbfFOSDadcjn+yiMmPcQ2vTL+xjfK9VQQoRzht0O6zl1S2pbHHuei0
lcEajQxlwspGfSRuO4dH/tgudPHRhHgY4n7/11qq9jURkUNBxlZwOgt1kbbotelewyUsS141JuTg
xnKeWANHhy35axjpAuBFWzh2nHkO6RClYIS85+NwPJBGmwFPtLDIDVGdQjJIyHOtlIr/MIU2VdQy
Zlv8BamgbABDcO3g0Q4h6uZLmEFuc6LQjWJCoJ82dZdDOKrekfyxiQ+6MvprreSjemHo76/ZRkNc
n+Tt6RsOAOudypROrJwUtM8kUoqhjdEAMjYOiF5yv5K9cYIovCmbaQepfCItKCNieYHenj74ujVj
CMJlVvIbdHMCcjvroTG8efnJtHWqjTIdHseWax8sdZsYKaz4FBSNFq3oMcXv1VeGd7t8aYjHS8v0
siuBuWPpyUVXwTPwPMguBzxobwWXZ+RLxptRG7ogSeR7O2Fwgbt0yhPmmFl99GUBVRMKGwf6+HI3
YATzjwTaZhbRvej0n0HZp3mG3M3In4cxhBnN9w2lMPz/qze6Ck3i7KpNVYK7JGOakxtgqjDrBaEY
ESycZcLH++KAQMrsTUJD9Sb4Kz+uMDO6z0OCyyKr5M4TQ5gy2SQEaCCGfNMkwEzQ9jyIEnVJVBmz
ko6nXJlGsnEPD6Wtu2caGcHTnfosBS9lX/9Rrhjvz4s99FyeMcIWP76d4AyTjJiY4kxacbqENFp1
j7f5nDV1eDi+ez67rjJLSEDI5nuk1tgksUygm2x/6IQXcPXliU/EXBK3/ApBqEKYHIBPrtT70jcm
ibpKXKCsgrsZqLa/CuASGYHAr2Ham2KJZvtg2F/2s+vtmwPofkQeho0Puj/SewWXr55tC4f8Lla8
JRHnAPTlCp9xQMFohynKqwZuC7V/tD/+0NJkhMh0R4A/t0M85FUOVMw8ZhdTiw6Tz4dVmvtAeeXG
EPKlb7RDrjLpkfbmfB5YfCWOTxFyPb7LmslLrjE4brS9SVTn8HAI6mzqTGZoW1H5MA9GjXS7TIn+
aFFI/LJZwefeFpQykzqvAH1bXrzP2CifgWfk0TNLstTGhcEmE0zkKdiOsb1hgtEYCrl2qXhTsulM
OCEFMNktFYtvnbWYR/MlbDjJq0yH1XD0xWp0j/VMG/JUqPXDOtaVUmRKgZqWMjG2ANHMiBk2T1MW
3Zf6DpqO83piTavRxDcEsQX/P8gQJu1m8DEG7O8BqOUiK4w4Iad7d6/i8aDYcNCHPk6W84E1n3Fd
pSfkI/cuW0tjKOljywUf4WZ2S6KGKIKV3oiVC01R3CJtu1iJB2K9yAoO9f/ejT4X+1AZcAyQ+Bnr
wQdNA+1ojpZOHWrtkWW6XxzbEJTKDMt7FZ5fTdp8of1GaIuEaSKa68rASYznc2kyjwvdmPKkfred
KXst+Dz0b1kvYurV2dAk+bLG4xBPLdRtQEd9qRRQ5sOHC9UorhoTRSGcBh9t90HdsX2+H3jpMMuC
VkcRDfYjJ87H/jejaJBlW+QptGpy18l1eeenNT/sAoCe7atGrOqp1e0EUWX+aW/MVZwKeOrt4YM0
YP58bDek/2ccHDu1vIWSiCU0AkGdvSeGFWsq9VXnk9t25aIsmLB086ocooEKUFVFi9FdNmYc9fUu
Metf9Bpmrl1zjbEF4aeoiPflZ1Uc3DdeMa0Z6qjOF3W5KeJBXh8knOr+6qajWEnckgRTV/9vGBxu
m3nan0bDL/dvadTkrt/N9bbQOHhCUvg1bSe1x754OlJI9BWM814TNAjgiduy4DlpJmuM1gmCNOXO
hgJ9ddNt7YWTS1O/LQ9XBRjHD1Dg/AFHZ0908w+Uuk5M+MC0+J8Q7O3pj7y69hekBzJ+LdQ5mxpn
RtpV3npBrpHNLuHKmXcCARC44k9j4HgbiVDQWiDdMiyu47NYpVlUJaaFeqjktdrjr12r7ySsJWLJ
xEZsdh3jfHBy4qdawrqRDr/n5lk2ks6olNld3lnDDKaPRdcrH6mJ/3GjI7+w4Yqb33fL+Wwzs5xr
W9Vx26gxf7RB88zUJyEPtqev5SFOgdTRzAA+Yb9dVNUJu1YNBx67L5QxrahnVVWYTVtZXV0tskE9
gFpROi+S1SggJ/VbWfglIKK5ivkCIhlNoCPmZhMztEOQgjfEYlPwIaBpDe/pk6ywFX9w1uXbaQtv
iiTRmOcyykecW1FCnGmapB/a6DVYQ8VotZsVhGwxj5VIFP1ZrTqK0QqVPOVv5OvAdET7O4I7otWa
LOIs1shk7UdWhaaR8g+5JXHk5BW+wtsBrFEBfYLXPwbbIHvUpYQNEY9/DprbV11QKnAIUy/WUy3c
+Ovpf7Eq0EIQDTm7GBJnfZhSWF/VLdV2lhH3hsjBSS801nq8TXH6EhFjXMPOTvz4nogKusjjO8cy
3qmnWYsHR3nhnnXdch6pBbhLaNcsLvqpC5gbPE8Nb+NaaYJVTM1PajHCsyiIr2FhmUvqkK4OomY5
qRYZh2kKE9ID05eY2U0Svsi+QHT8RMiWcQvowqe+AfROb5ryCBxxem1awoQ5YXRfx0ryGWzuWmXw
XeFWmYeV6qADeygZJo36ToNS5spRg8tO5b5TZ0U7aPF4E4E61QVr9iwBmy9/Q4H/OGArmM4XABd8
vNbRJ8UEX+vgRGuzfAAMrA2xXJkNuLkvIPVpLtQALabVlHe70N8JNXGU1mTL5A2qBsvHXxeMDVOu
Z6ofAinufZg63G+6IEG/R2eSkn8uGrYDwqSYexcs9yC5DhgQE5Cb7YRe3cEEbC7MdItsca2ZT4tH
gy8Q/zTRbMgk3Q3ctLbrqKJ6fMS24HghrkXYJdpLgxFB5WDDiLpOxv5bXOrflVuvgC6qa7pZXn4F
dQ3041fWYlgdSGTCFT6l8nl2tiDSkqfsX20o1ESzuoBwQmQTkK2QououAjh4a6TKNcqRL74CImy9
2oFoD/RXXkRSl5uphE0d34QyiZS4/yB6skoJIipfEGZm2pw0HEawZfuFZtX0N8hniZJjh3SrFH2L
FJCzffialjCk7deLC4Du1kPT3EXVJ/9jLbmfUyTK06qp+YsIipOnqt2MrLH9b/ZHiqUBXoamuKvp
SOEy9U0Vi3QwzuFAODXsj3UxV6IrU97ZGxdMDu4W/E7nALiVlLnIBMPMpnyRjBB/+j+bVy+cJN3F
2oYKAV7meQeMfqCiFp6dm3LmoeWhcPZyUtdwlGgd7IvLTxHLeKuLgbVAyw3YumwZ54JTyNh33lqO
hjRRjuLTC8orc42x3+qenQqBp0ifR5erCSrRmKj8sR7rrGKBpMr5RDTHFsqKh5PUH4TjW19brt/l
pyAZ45Q+e2OrBwA8U7GTSJyV6hM+THNLL+r0vkzW18ZSfJklm3Q6OrQbhoUbSv3YXIJ6f3s0hF/i
NwIkNzPa1LSDJ6oWRIUnxIkCQBg7QgUVlflk5PYzrQ/I961yO224qzgl7pS2a5HQQ2ES8ftzcxfj
JxsRopEmPcKoTqZbBKZ7T45XFfHHEMetmMy7/ZR7U6Yi2YJFZJoEG4ZKYRVhwAFJNZ82QZX0jwLz
VX63kV5VP0wZRQe4SYgy7LnbT7YpRFDnWQ6y34FlJPx2iC2g6LHgumBu4sSaemN55YuDkWYa2wzx
hj+4+wcHDGV1F5UybB36isoVnTJWBEfZsCV6kfCRMoI/GSnsZuO3a3By2zzE2R9Ybyl5dqPfXIzJ
nvbkMDZh30ZznSKxV1w+sZ9P4rV1chIEgRwsEEftcmlcp67Bc3Zx5eOkbdrqSPwqLWlW8gbZoEi3
PAZ6TwJBKHbw6312BtKS4V+9QbK/J4Jrdqp9ytVqF3myeI4mSYOSYpifZkx/qgemcvUc64Cenyyh
7wjjdLVc4iQA2L46IkgaNQg10T0HxMwblt3gh2YO9dmCE7uImLwPgNA9ZT5JzBOwhGrm/NAuZ7Fj
KV2rTKNfD+zMhPQVX0b1bWw39X9mc8ayXqTF7NtPNtsWCkE2F+4580UmpZvbcwfu0KygEZIcjdr4
vBJw5146+csfrpFWu2dbpkPqXlkzikIxsCcpcFLWVs+zfNWOrydZdDTfBABeEuVdG+u0NWNL4ptU
wHOX08xVydNLv+izhr5Nw5bngmJq2myZUEXVjiMd/SCHx0CXw7JXlxFtz1k6da3eejoJeTLDLzhQ
PQc2ImLFVMS6Hj3PIcTQYtsjnX2uvnPs2VW3NDNY4Hiyd84SZtLIK0nByDuR6TBsZud2J4S/aEXl
8cKl22L4C0wxkPrwIl5N7UmERmZxHxNNidBpYTkIkv2jiKbQkm5cCct14xrkcB6Pd7NjraT9wdQ/
EPZFw0M5Ibn4cyGhANa1y4CAJEITG3tjLT4rUGHb5PIGTWZ5sIpQrSUWSf7fSoAlpGyFbLtRYiNN
TonjOvIPBDMYYQuSbi9BrOW8OHuGFQbfG11+M0uMvx4XRYwgAYwa9eLENtQ3RYuXqrBiJR9JPssT
090da+qRTBDpUYXaXNjbXcZmmUujcxX8Qj8iMPNYZy1mErLXAVrZvesJuGYScdR8VfbT5fLVAGnk
uxO0+4Rk8nFSbvCM+WY4Tay1wOy4oeuRi+yYg9+2526WA92kYv+za0abkQbTu7tcF9HG9AGwIArq
9oefO2KMEr/aALEpHrduk4aorH/oxY7HxUYVzvwdg2K7L3RmiFUU+4d1MJet2U+/QuhBvcYpG61Q
cuGDIbSVPxluUqHR6lKjpoT3pCG8LpCPFd9wuuUqX0dYNlgKaFlQ9yUE0sVmUCWYVlLIC5JGvSYM
Qvv7HrlAeH/FBF+Y+a2QfzlbMNOdqD/UEX2RI0FBZfpmVESBNRo8utrpBRzilocK339IlP6gMicy
I34R+YCV+LyvvisuJQbK3ilTG8qfkRgbOGqhHzV+rmPrUGLvB59XakddcOXhQkl68EoHn3anDDZs
GiU9vSQz9kxk6kx5imYs3A9LBknyEz+zE+trFhhzeJrDCn8ToywFP3xMOgGyRhNLnKk2MqxSUTLw
1KzXBQ9Ts2gUffgD3ATHfv6+G1blFkZlDRi27R1lDggjnRSWqnGZNVPYQR1vAdVy/3hIiweNlSGa
RdwklPMZyZPM1YTb6/9BYH0te/8hURO90s9DytZZyuoScmAEtZ7BLgmBzrTetiTXSu+Ic6YgzmRm
5CXAMj++7YRU9dZI3yndKr3mWk4JEXtSUnb+4/OmhrH0WJUmLfc13EZV9wjGt23p244Wj6EZA3kA
aDQ3W4GXRU512LRUCiGKLg8GTWKqvL8hQCexFru7f0XVg6Gg4AaLohxLEYNY/SF/FigroaTaKnz0
+eNQxIU9Avs1qq+cHJE4GBOeUA3ntVjNVNjRyDhsD7lHL2gYzirAnWfMjBfK6D8gDNYuErtzlvBg
rLp9Ob+Sgf9ShQBgyjAbPyL4cI4U5IhmGvi+UgLluJTVlDv9Lw30e4WeHvT8MHTAgjdsHHVjGinU
ObcKCJzW4MZf+WmooNiIV+vka6nhfCro2mhG+Ww5+FT2LtDM8xkd3dRBRjO0FvTzClvyPInZbYXv
qRjh2qYG6aLA4rhweuh2EDO3YRvwyvP/Hc6NyVDG84SKxWA0WJa51R5jkuc5mVA5f3at3oYfzWji
wC4+Vw1LMWtCnXIUgWOaYGzJd3XDo9CDal6jUUtDWEwkR965g/8QZTj+ckOGaexawsGH/DPFIwY2
yy7R4gpzL1xTyKeIhm6o/wsPCTbJTgAArvRTJ4wDQ+T8VKPpugRTUJt9Vd24CzAbByGDjqlmTnx0
leJFQEjS0IO19nAPaL1LDknWXK5e0XdDyImzoBiXXCV4rmY5lIXk5cziqQHWoMvzdnLDdr4lFXXU
wugRDGqfSQmRE1dVBATX7CEylz1e92hXrFe+H24TD9zspf3TkXUIwU5Q4JbLKzmj9Xk4ro5E+2BF
nHghsat/wlH/IFsb3ih3qVMgZ+mHMBPpe3ZJyAf1ynGbfDI9LuAf2hPM8YjUv/YMh6+bzho18ZS7
wDgNQr89ut3QAEKhhn8CB7lsqlKRgBZClVAaw2UFLZiTdaRmtpZh9xFpiQi/47JoN0zYiz6Sbg8a
OnSG0gkWrasUuh4GnnloWzdufz4tTXcvVdNhFBI26+VSSTxFoE5pDEm5GidTkNlnMIPDxhek+jG3
m+L/3VF/BnXIoH05Vnec4bHqH/qORETfL013g5zayDXfHpKNS9d3gKzOCliks+pVeFoKA5DgJ2g1
zoV0QejbrlvLUmgsL+x/PcxT5ANXsjos/8dsZ4ytXof2B+qL13PladgMTDZx43cAx6m5DvSeYK5v
0BoYIbaP39aeMz9hO1dZnRvqfqaMk2lutGsvpE3a/3PQvdo6zvVDlDPMaNJCVKRy9coswIRVnxay
PehrJ3V34Q2Q4CibmGtuqYA6kMOloyVKFl525hsnKhAwvsc2DuiosOrOfpSxqOtzSlxQ7KnzS2te
um02/JAly6m/SyNTNs52GNdfLSkz8drsCVqKqpKG/tMEiE6tSudLIksqWXJMOAR0yuDJzSsDRgq/
6rxR4J1fJUtGUxXq+5M6xZMVMCaanynNsEyLEqL9ubpiBMvRL/dUi2gOi77cY9n05W47Zg82lI/C
wqgKoPXpnng+fuMm3aXYaKI2lDZyMGgFBcbd7bz7c6uWmLZHJUZE6XViJJlzDQbtY0bcKc1C9FaI
hDJ7dBjr0qGz9YhOOODPEXPIP9AfJalqsqiFdkY9knFrE14+yjXvuglM3DrL2rDLOxJXZ5XPd/Du
Qk9BP2vZvHn3Sem2w+UARaccUn/EwqCspg6yx29KqGzcmX69Vn32tNX7nTnJ3fBznexHxFew5MbO
HDTvEgddAVHM0oDMg704oWmr2JGQAQ6oZH4VtU8Hhl58nh+lVzCR498hV82xTUyznkSjs3I2bW2T
YYUmUmdqApZ2uywFlgaamz7lS9mk5pjw5UJTM+F/dDbPXPrT9T+RtZfdWBxbz/ZkfjBnYZxYWGdx
g0WGnt8XanTv3sQFSV0E3E2zMfFK/rWBX+CdAaZGJ/CtWLu8845wyQp2z3w++AZVUNy1XSUTt44e
v26UTk4NIr4nSE1jRJySWpwSb3eRjW3RKubBxHzHeMdPaBIZSFDDdHCLK/09JywzQwABKvwyHyIW
zO4xkogLxMUmyopMr8iflhGOE6nJG4OcQblmC4LdRINltBQYySDPDm8HJ3GmXwddv3XvRUle+6x1
FvASRaxG9U3epUMWVCXapqZcr9qHwq0HUH7cvD+pjNTLahfKO4Jw7raKnPqzunYRst/LtTX+KEGO
MTKvM9gCjWhUOFRWscHKY7XLso0njKcsC4BsCdnqKiFzSgKamFt2fG1RyzHdg7Qxr9pOz+v0o5FY
vtb4/OjSdH2jxQgQpT0DPFFlvbuHKndZ6rsVvuCR//lAnDvxbWxzOdWtG2HFeWPUhQ/HG1xyKBVV
ZPb3Gi/H0tX7XllpveCrlhDJJbK8Z9NBo97MvU5j4ldLWzQypiBmpIs9DJNooNqGODqnRL/oEPOj
yVHV0q21HZkMS95sEmnWBrSaXRNAqdX7ZbIljmIr34kb7mYqBgapce5SorvEdrLrRBsN4F16lsLT
eh6LvyXhWYZt3rnZB3FutUzTzG86XlHm/WufxxGDKk0RKzUTu7FHKglrnCoskOXguB/7XcQg2K1g
TtaHhNOj9VAXqA+UbOcaLonSUBfmY5Kpm9UZxILPNlUWU6lLwC2aGleXj7HOQfCkdm6j+Pnr/Pdh
0OQMt+fJzUP/Q3JDguiMmQbo8w3wc5ZmBdgoIlZx99cX+SuuPtJRrMSI2/dLmB9UOXKF/owdxT9d
2U7FxenCGtevRkGvqu6dTTZf+ao8bQbgaJuCcueVaIUEMssghdL87aYgZVJqZZFboMyx5YqDFhfg
W6D/vIHYtroitAB5HCd3uPlubXiTOTIaZScqsdFKbRA5y/xdrgaaS8vUkkguIHyw+zdvjcQR2Smg
zKjDUSCwpHC1WzxVxur+IU59ThZ6RgNfY5xhTx9uoGOCvcg95K7S31cQD6hbT2wNdZ7hvyGJejmA
pUgDkrxGIWfYjPnN2dcCwrhtprQZh4zsWJwTUErGLC8VxM23u2hRSYHJ21LbsUk1u+EXnCHUEWc6
S7GhWrnm4S0bEIWvjKvuSQNBUr/yFVl9i1p/67x5eSsUKn2P3hI5P9PQDMCtINqxshGrZnzfiAJD
MBCWZFbnp3jX9tsx+efxPGpCeIftGygO46Gn9KWNzNDXiZnkPmvLlvlIHCarvlh2aZPDQvtOdvAp
1meLimG19vGX014110/cXwXagaYmfGzcXGTR7U4ij2zGaPVq0O1nHPd0XMFyNgCYw3m2TcPLgwmE
sbgC2NwiwakFmhUKhfThkRL2CYIUOrfHndMQt5LWb3R52tDgoNj90aH5texVdnQC9qfuQhnoeJTW
WuurKldt2Lf9hpkhpaQElN/6ftTaWVZTfmbMJIscbNUSHmQ8DyBAYE5Rz19UZwexMBqdy0G04JBd
IfJ5NmjslPEV7wvLf+xL/X7zJM9gJPeie4MWx5g+f+0ghZA8KKugQ935/LrexEkRzICfeXkvQ8Yu
duSOHyTv4f7e8ohRb4nFI6Ls5oQ/STwRvC9bWIq1PCH36UXH00L53mpKk4UIOsEMmUTFOlXCiWuy
4dG+w4FkbjmnoUVL/19ybk4c6djcuGTY6tEYRzP7ftOBwgZdpPmmwh9lQDV/zw/rA7Z/Wrnk4d8L
ubccWfg2IT4r7hk1+Jmqx0cU2Pujse/t9fbFSWGXhJNn4i0RQEa3g2pWhrFOJJeeLDvqW0D06pNh
8YuTf+M4/gGPP5Pgj3i945ReCjKEOU5mQeHcsLRtsQWteMgdd68l4DBFqgb9l7ioKdOuMWBs/L7g
8DTft8hr3FZyDntTFUc4YaMnETvKdarNKS+uWkjlj5nQtktUyeR1J05c+lkvf0feox1Pyy8HdjBG
JVutwgs9BHeEWz73xaGXfShn+JGrhPuANRj+wtlsBneeqQioGgX6cANpMZQAKmMTr5K0/cPyz4va
1wVOLsv976FO/xqZx76cjMp5JjIvrCUPXn8quf0auS1ooiI/3mg2tYjAgPjGdTS9B4lNGyKQZJTr
eExYooMSK+fnvDYzKvLj9uXJS2aRWRkAILBMN7CV5dvzJpZ8lVFSH/JeDDj3xJ3YEPQI3ybSyTVT
Jj1wXAVKKZsUPrGhFXKsQETXOppGo6QfSSq1/k+tZekN0o+FpIUThHpsCz+eVvqBzTF8R4mHPL1t
vHNZdGD/BfMxkTIY2Vw70rM9uxvkTAMuDKkvPSau7tRanQsNCpVr7PSFd+spEcmj12t9auvlaAnY
dVQVnylPjo/AzF5PNv/R1pB0OuLF/4HLGRuL6wxqA18ZnpLPP3m3TObNvL2gjiugxkxjQwirwzN2
uyUFvVzdbBpod8gsr5QCm5MdUlVsPNX47j/+OdmjGNekgfUWWByW8QO/aM+gWKNaXTBHvAQlqhcx
tULyipXK4Z48jdL0FFJZyXiwPWmSEg==
`protect end_protected
