`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iEjoYdpoxcGKWZRsp4oxv+EZEzUSeeVTTkaAPRciDJnSfbEPLLKYk8WjFSfy5JIAkkCfE3q0nnVh
qprJuZXAhg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e9ONTVGwRJLTG237UzoAJdABQ5rkM6DnHXF/sF1/uVdMNCBT3fG0w+FoDhz8kXvk6j1iqmQ1uNA9
MK3DBbhknUW2va8MH0azAZdGR6GBdKzGZYE8QuUtH6j5P9PkRg4SZTnRUtqO2jJ8RZLOqd+teMAJ
E6o8SRMPuN9nafQBGnI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S88fbr3xQzQUmg9JRSN/GAfY/ZzDfycX8xGttAB4ljVrK+/Ud2wPf2T8zdM9B+9tK6YnyyKTucss
I0M7aYVXOoOJ619pvkbCvMkvYup1ThvrvX2r1cAwS+XWnXhhm1JU8GTYUnkF4TqjhaH76Yh5u/EJ
DkQ8dkPQEL8szNDBY37WanHciweZteIA2EQ4bs3Ao8G1B1hOKp3n6vnSZxJXhpdHcqkaCUufdqaM
FrinxwWhd2b8vF7Oemr3OSlqM845sfCrMN7jxAAgHLAM0MSMgfKTq4o8CRsTHWQQzAOPoqsx4fzF
mp1LX8/oirmCsufy9CIJjtJkQ5LMad2v2GOxng==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C3UZmTnXNO2JOGNm/uXG4U8HlhAkjOphRlJCOT90GxGNHlPsgnu+YFgyMxXFTOuWMzkcEiU3Hua2
KsBVrQZL/9/nADC8Bse8IldxE8W/BOHRy1TparHAlHZ8f7botWVRTz8IoKsY6ckC7flbSTrOvlyz
+5nXc2aXR+lsQkX6n60=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sRP5Gn9NwCjZeAz8hSSnN0il59CdKNjwYzXW+sllZnVXN/N5yMoHSeI89GYIqBSGSsb21UVo80nC
dBxojivyuUfqpZS+t8++R4eRbffR31bBUrrSVg5OosCxPxSCHv5hLr7xlyVNtUmQRka6Y8Wnyy28
blH9if9JaVp2t7EInlr0a+t8wf9k5dP5A+bQyuu5Kp4nDwYAhs959ckVmufTJxVslYSH8VAMtrma
FNvPsmO3pTxY7bZ/PEIDLrFc0xA0mvB2Un0+Z8TOrxywRFfV7kMy4JyJOJ3WcAqeFWr4la5LuoH9
T2OLtZeG7TTN6g/8bQwzuQY2sSWtxugM04q/Jw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CTYJN3IGTSMmDt4BcedvsCRhsSnxHT0LScK1/qkByuKrhygZj+r7nAppYsaK2eQJyT5AZNIKYyYD
PwobzSlRvdtK+Ju2XN41o4Gj3J73RzyJgni8RHg9cUcf6lZfEDC0NJesqtbaVfEUy+LRJkpkmdWU
GLgqGSDsnf7fw8RjZ+9nxPuUCJgbOp6zwafzrF4VL7aYffqyx/M7Z8fxyq17ga7TU/prOzR35ZIk
uh3XOxTHUbGjUroCj3VA6LZo2TTNBh3OQZBRdL6lGNwRqc3B+I2bfUE4RotHIOs8kqNPu5I0o5CB
G6PFbQ/NHr/rSrdVyogIDq+TPL62jsSQ/f/twA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 115888)
`protect data_block
+W3fXb7xlQiLxlTFROgPorxsH7n5RnUufc8aCIi8FkOG334azkne1vNsBGoZ/rzuCf3KdLB6LF2j
xGSfo+XJbmpKgjIOvSi9/RirhJex2TDreZ3OwbVT82thHSZY7+vu3coShRSkAMe5Sefm6Xv4hnr/
jt4YVqgaDIJvd7OD8xSoNzG3pZzRS+qbT1Gphob9vplCUN9KgdKTDY29HnCyaA3PWLLBOND5Tidh
YvLzlEUz9LmNQuedp8KcXeJAe8IWrMxXK+hxuMUCR6admVfQi+3cNTqyJZUaXGfoTNXKS/ZbGgcf
6aDOiM+Ot0BqGz6ogMVUexxBP+/DOnn4C8/doinEIwxiH2sVa1lmzxOScoqK82qr1iS1xnWnAWng
QAGujmMJZxM6aciGpxj2yZRpJAAZtU4Fp+YWf09tERLTjyhK0P9Xdt+DFk1iwdUXolqkW/G1PEEw
oshGVgnu+9HGfMRN3uG2vOB0raxqH25h/0vKrKyzIau9D6lURS8c18shUJTxJhw33MjE42GdSXUW
scErgzFNr62r2rzo9P0ydChjRJL4mN+d0Lhns/OH+8DyoLYxCJ7qWeYFduTADo9a9yQTN7Rs3qDG
Zy8AWLvV4HYySTtyYzWTFjxgAHKxJsWiASUXo8FdRAFkbBcXbpEykQON8y/mMccd7eAjgJ0z1NKB
ZP04GrsVd4WvWpGAWxST6Xa7B8ocwO4AyEusP3B7aPK8XXixoN6GAuZZ6CgL52FfPNrkWAPVLNam
lWZ+3qblXsl6+wGQGCBaS569y3PDxQHWWWX0c/nav84BPXCuxWIYdSCNX3hc4Z1uf/tcI6ecIY/N
XZUogTuX9BKErii4HjfJmUIrcMsv2+aoGHUgY1StP8QvVC8ONXdIXpEjvg4pC/FJjwWxpVls+KTX
K3+hJJo9O6HaIRgKP/dbMGVS61Tb1RG2X+Z4v72x+KXoxQ8S7p+T3mI/+g7mswUpmLfM74f3Pw3q
n+fpE3dCEzzGT00SQUho9r3nylmlYbmemAHmTyVXJbXHurCZd7Zv4RAD5rZUSv8I8Jge1w2Ocgpy
pltYDlPZEgADotuF5tzb4q4J77jMfBM03wLYG14MobKWNKjJkvxdaSZgrD7lUvXYaDRSub/YhISW
uQRQfEpWN9KaIW7eLcbtzrPla8YQyuXhlF5tRmZs4uXICzpYc/1r80NPFeasG7SYstZ5/RKbQMDb
7YqGeYwQz5vfBK24A3XGYu06eq28ZvtA5akOvkHFlD7Ep8ryo6o68FfO4i0fcd5ZmbTVkScgrMko
e2qZap1KR8ARceuIuVgqCpBqt0Qcktg7ySQjhiunHQR8jFtRJAnp703Py0xKkwykXU/IVpzDyifF
EtCH5OPMgxLVNGCv2HqqSMwXI58FzdjMhK4LPxG5DPU0nsDe3HY72ArQYVE1tTbvzfH+r64fYa6W
lPApFQCne6S1EamYE0+zFNv7iOwxRAMWTFRPHuYjuMdTSUAG9PSG1ntE9j2t29hyq8c2TAOohqX/
mPyBB0MRTbpr3E/DNOKS+Fq6yeMSMiWUpO3fJ0v5XKm2Yn4MX67bwMvEReT6A3x9GQH46V04EaZf
3yxJxL4VJasT9l1PNXfUyflWrN4zRYs7PUhk/JD8+9HVo2uStAEgikX9UtW9G5rYLT/HqkIzZq1E
JAHJx2ut7aDqAdGexXJJSnSKy5DMrDPBtdyMuV/szb13fQneBhaYjcb0VT1A9FUFF5zNT1qXSTkY
qKvyzH1EdzzbcNeDZrVy8jrvEGgPLrRy5H2jrSZtMS/0MSr9hglPFv1czSXVfmIHX8shdct1Q4b2
XwH1BhCw6qRBNeS1iWV0j0JS4w4FVYmkbo5TDPRcl2IEuUmy5KQIWXTp8Su/8qQk9Y4RPn3Jv6up
txG+YGsf90dGO0AqgSgQRQyBvQ4ORqKfJDihun6fRcNVqiHwir5xh5RzJ4AiZJuHQRxgWeHeF4jW
K3C2h6/CDWAvjsQIV2tJFDW/2j+OkWAjy+rQas+3phBQxL1AfCtT8LqEL7tKdCBY6LS6pISuoVMQ
TmYPfuCqbtgzKo07lodGQwrQw9KivNQXhO6dHP6/Q1oFFQTdYdVV0P2Oj7Yhk9xi9UKE1DSbP1QQ
19rotodGQVIn+N9xKv84JN7ujbo+QYs9cEfRLUn6p7mh8FmiXgU9O/Y+PEWtByMkAGycBsjWBG10
o1GxZN2Kk7oTFDftcYFuCpW6B0cxUNj29YxpoWLWciVIHsywPFMiZ0eWOJ5+prFM51vLsQulMfhI
G0fD97xxqA/BGxxr1CZYvqCrKAf9cWAQwkiQ89rF2UOq30P1uJZs2I3NekfaDus5SdizvbYNQblf
tcbUDI5bJe0JcxMiRKSJzPQBaBgDzAd+7mIV9C7rVEGi64KMjH7foGKLRyM6NtJeMYRCPnWcKioB
FEAOBiZmGAhVWZSK3p/n/RrmRk1WC2OBFftow5TJSDOXmFVXsNgE6vJTJLCTpZKaIWIAXSQE2+gP
0F6OrE0HMugPDfzcskTq02Cu3QjOO69BLsSeg6R23kQ05p6d3WONiUH2GFfh3GtP5wtDH2WqPyU+
qMl1AtTEfdlmdRnIhuJ4/cs/ovOOUWSYC3N7TUunN4PqmDybbxM1+KzjQa4HNe1g4JLE1/1k9Oq1
MXI5NWHaHfT+lryfQWioRf5x84X/dXWwJlfeYJ0xBW+SmMEtWoXszDySbBY0pFRZno+gSzqUw2O1
j7/B/5CUnH1fYjpHDkbEHAO9wNGLOlSvNoSH23fhIUmDO4whZ+kBSskDKWB148cbi1cl3XJlVYTR
EVQ17GpNXHZGwgkYynqFocPuAnuU2MRW7puzEtOMQu576XOfY5ewl6fIbK03QJdYeMF1TJDcGJJl
XGgfAGiGwFotLQWsEF7KueNtZCu6sq/EcoiaDhi39sE8LZkJAKPx09lwZZjA52FNpePpmzSej1TX
e9MjO1KeIxnmrVbGCstJtwMmzA54wW3Jg+Som+lvbYYnTr+3okIeV32NF0VPyr+gEYwfr3necfOq
YbRs0vDqkzE6ncbbtGBC+v26NqEHVrkfdNMO9np0ZqkzrElNI6FHq4VU6W/JP3suar9C/V7WYZq+
fpF7VOEFQ67NR/57jLndAIm55oyNmG2Mg9YzSa7oI3zR3pE/p6BUo+MobK9V/RIRk9RFWqzzMxvl
/mufo4sFvNa517MXqJ4a0+CHqEEsBtii/ps5xz5CTTF5SjQAdzSmkBG0s9uwXXEG2XIOnMq/MLQr
F+UzlwRcdb2ajvovuT3KUALr9W3EzB5w0Ca/q9DJOTdEfZiwWX3FXdUHP+f59G5XDxXv7Lx3iAGQ
oC7w/EJvmxu9J1laakdPUZN6zdc1H0hO0fl4lPNu7pCklHrHeFnRPSJp4zoLWIcD+CfWNrgOa8fY
ixdFc20rRioQxMo8WJe9uWf3IodFHrDEYuQyNuaLieo/V2PCALkULn/45uh5CPALy764rGDPMRQ/
H0jZfn7qFR3W6TwVpZh4zHTH1EJTC+5JwZJ7eq9rTyPyHAcl5F8MG2tOIuUtnvsqWPx/gDI501+c
Bw0vUXn6oYB+/iY+inE0kgOPXp/jry4skeaREZefZFR8YFQpV9q6slcTDo13BTV6+17A0qhzMzZN
hKkSThuH94v75Cnx1+/mAT73+cdXYhYdOOrXbLjg+j1j+5kBG3ZfdbK9y/oZw+WMALGCv2b/EuCn
7ASIskpvKu2KILT1SoEKryQp3Jp87vwrnYYArQGVN5IXTwB+YaliSPGVbqnVEAYFN6lJKfPGoES+
aWd2NbbX7qhA2Ws1P24245RHfvBqT8s4aUam0LbbKLLXHAHRQ9gp7BOr/0cUFUmvrcOBGVxO4aPh
ucJ96uQg5h1HvyrB3Fnl5/EQoOVgr172MhU1G/cycGZkSWNiLznAovpBoWW1M+3VjTy9LI23xw0N
m8feBO8QVWVQd8/M2H7KzVj/FkHCGw3/nQyVCk5+LO0/7mDAnXKihOC4Y0ueQbJhC2LiYZYS4R4R
ZRWsfmk8tvBopZBqLtUzOPLn+VXRvk0t1cowTQBPE+xzeCTqXrDCYKE3o6u1qkJWskimC55PG1n7
V43RFHO4NbhTHKZdYNBKhlEIahNqwIyPRl/yA8ysXtuFVCnnsS+Jj4JTa1wloU5fxnHsJ9Q43IUQ
b91ZrwQIwOXqzORIjxI3+si7j67Gvsulf5TCFXvVlN5VuT49Acb/iMjmUwG3uc6iDpWaxpjYakkp
mDyVZF4ucSfxYZWfZQ1mN0mMd2PFwK2CiCTHdNrmsklw16IQo0TB9vizO0nN/vNLsKfjjci/8ayQ
RZzR+yQJbeCET/7iWyw/ykpVfbEjiwAQ+QNmw2lUi62d7qp11Jn8xULWizFw/pZTRlC3GUkwo7hg
/KyH2Okv7s1J9uO+rUmWDjn9nhqJwqIJyGvDt59s4TRvTXJgiT6Gk0VB1G0Xn/HLDXV1Mf/8/LZI
M1rMdzKSQvKWsyNorfc2KETz+yilgo2siMbPXTqmHTt9jYC6cOPSYHcTdG8uSaQ9/DViFmgde7i5
PXGGogJsIHI6HJ7Zpk6yuVftCHsHINsPLlK+EhyFlDBoTlG1ONFQduuKbscrgIPNYMwI8WJWj/0K
SjwKpX30jsJZDCkCh+zhizoEdhDSxzEao/wudXLO66nVnAVHB9wMAnsuZnQEkVvySx4YUJaXHimQ
hv1GfQgStjR4dDvqn9jVPpv2W5B82JgOTeBncFl3uCJ9zxgJuWT2+wE8bICZJ/YHKq4nSQXAvxbK
MeGxlQ8JVYqK2aFGV6nJDrWIITl5k1mYjpCtEzBQrwT87VQrK7TYdeDBF4soEOJCEuycis310YX3
Goli7LvD5tX8ZOMcRUHIsD3Y4ioSClzeijCzoLKkTBK7EoGxBJh6v9/InnWf+RxEePtcjEOhLrFs
iUDGG5f9EGaF2w0PiYMqOCEiiHLW4Pgrr7lmSzv4tlFjCrHkgcqfI49LPcVpZLoRs8+ZOqz0kgLc
VMCzcci0HBAEsoWifqJRJ01njUIS/gwWJTwOXsoL8bSqaynCfksYPVnb9IHnRY8RuWkadBPVB5ln
d+qaj3hZkhKctyIW6I3ERLAdMe9hHi6N0i2J9KA6/2wZpybMJuEPrOCsqRdRqXv4xIu2ZuyXvi0M
HVGuq5b4bx7C7xj2T7QCeJrlnbsrWQGpVLqVf7goFjwGoxrV8CBna6aKEdr6DL9zQsp63mB1J4Ma
rY1jRlR5UVUGX8sS9atNrsSBszkzNg1jcUGxJ2F9Vu6neZbA8siDuP47LKgQ/iYN6Yhb+J6M2iqi
0WRC71QUUtRvdDVNNSLK+2zs8csXmGtW5JcGUeX3YJ5xViXXbreJj/45fe3Hrj4E7wG/+d87QccO
hW40rc7HN0l2MUkufhI1Sn4SeZzrLJAmeSFBRyK/TbbPdzDH4ILRzW1gW537kfynXd8DCX56MWBE
scJy2YIzsUb2YpR1xm71vJ8Ex5q8B/z7rAzZVsw39NpuxQ4KFgsfve5F5WoMMxqAfTYKGuvZ6ngI
SM555uyN1Q8KqQ+JxUWMz3IpD6tgEmw0boCu4C2f/bAJFXfO5yRRtdlkE/cQcDPr4paESWPbo78d
qDU3O6jNHsK6ZEmj/iZYohmWMbl67qq589nLIrm3i+EU+YIXlyX+cB2/3mzKy0UMlfHDc7KQysJX
dRynZfuoPJ8JX53C9Tgh9LQkGwS8OUXm4NP0In/jjHY3E8C3WY5Ym37sfr/GN2tbPOpb3TeJtb4V
HlQNFn3UboQJn5ei/ibhHMtudvc8OZghN6p+iCjNagNEgwjyUhI8vSTtlFqUqMtbjA2KSFV/hmjx
j8iHIGMwIBFCORuX9Gg1n69alL44Q8kgs14OnnAX7KJOrxBNmpcCFyY8GnuYiZIozyGSbkIocIi8
U05s28/gT9L86jvdfZSvltF5t27w3Z1jpw9fBZzp5uXPiKy8Fn/Ii9h+qEf6Q3toPRqcd7rnmygr
Oo396XvkeEK/QKwFV0ND2ct4hkUtstCYLwFLYfo9qp90TWk8oRgxZLe7/nzRUX/KcsGeYJdwDWCu
mmAyQ+grABcLULNqMxSfyv6T+BUfaOKILXatsVP3hiTwsRNY3QkaTY7NmnLzkaQo1Di/aAXT+JSE
bgp2Bxd5wanbkaJMYAPtNvY9M+bzCy5IYukeLV5NJYBEorOUuBnQSfP42cE1LddAt/EANM8HEv57
s+AkweQAotyFeeF8y5h/lwvoyvt4PTc22jjdzLMcyaCLayfJS8iwJ4BScF+C6fwxTc1l2HQUsA4A
EAi9fAo32REDrSi9bffWDOQoc/mVTeU+pjU7OfHq4O5mwNmndHpCRHWM67VA20xa0/VrNiIAkuh6
RyM7SduT5TLKeDhYcW4JgFl7qRCkno4xpvGGPRSDKXCVNCOgRcQVLHuJ2bFdVs8xrScKGMMdGfAQ
AAkJG9G5xzFbeB7jaZnzHffvTxix/QOqU82o+0n8fPRmx8txJNWcx9nNoKORwlo1ix5QUhzoq7OO
AFfPXPUOy1RYrBx+jQEY+dyY5JriQ/Mkh9e1hwH8O6HxdXmAcM1JIYM0EfS9LkC1tJ0T2WCNTZDU
sxj3YK1bsJdyFM2UD3eZ1PNe4EcorzxmuOtsZF3hU6uJ3O/TPGlyBtrAt849jnL6K6BMjp7PEQr4
CgvOUiegGNaMjhjSTua/zhwDZ7MqValRKdos5qViQ3O2N/nH81UxKCAgi1eZepbiP3WJi0Qg4/rV
yQeemmCdAtXj2QOgJjRvIF/wxjOmV+R5FBThAxN+JPaoXgGm6ElW7anOaf2xV5YrhCKWckRNO/yn
clnOrDz0edYEan9M4JgzDd+wdU2PFSQH29uA1m7KYE2TxQmk55jvmJMxgDSc+6qufM0+9qHG0ReW
VSvrGW9kw+XdyVVuDSdRTmG0cwsqTe8u/DkW50JS279Zdyug683VBruu6pc3sTifGr0E+Kec7Z9t
D0MG2QM3vQlfxKYYaSwsYauAXxrP6F6MOiAGAGnthPGKmVlCOKdt2kpW98q62MR/cwXElcFp+Bmy
tRguzXFf4FwOB/XElyK97SCGcXIMlOIrIYMFI8KQbDSVeXWaA2DIzc0Lj9XpC0Mn14zmMy8AjKoH
TcCpUMPgI7cM6bfoQDd1aLDlu0o8fi6IUaFoOczonbSfd1vFsUdt86VhiEI2g0REdRelKGVjDGzE
TsOT9UmDfy5wWyJ3xsUh/q5MOp4TmeQTXlwGGZWXZkk5fJVAdtgY8Ofdh78vzqmoyl4o2bP6Rb7g
VZFrKrvpRJKShF2kMg9lX3AVJSqGJZ50NOUI6sjO3HoE676Klone76ba+hnlT4eA7/91tv1BiaKs
QNMgWuCxL/Igc/JVH6jyDxjrLtr49WsRTTIGThiokT56CT4aQ5qxkB29WQcikcDduWHBxj2NLLZf
B3TUaqyzjXn3cWRyiJ0kbNPyNtq0MyHkhLs2KS1QLZKNufRfIKRA42qisoN4wmjGxjkuBDP7Ysj0
KZFn9MtHAMnrwrkj3avx5nSQnwU5ca8W/ehOC47CBPXnnAievldX4Lj0fYbISrPCjOMAOZRVSvig
LYDARUUZRQRLKQxomQKW7J20pcR2xjzy4U6jTxzszxEE19Hbi6y4EuyFn/1XnG/bvRTrVmcltdG4
Sfg7Rit/+NsMItOKMdPH7vwqXJ2dEjHwpGs3sKxPpfKNngK2eVzmohwatMID4WfKBh0t0kobavcF
X4Qyp9wNeQi7T1bqDp9ZTmeya0xUWwFVChaT8ClR+gVKjVlXWMJQ6tkrL7rhx1IkMuN6VWU9vzhH
+LOmsLQ+w9iAxK3gAIlLS64IG2FvQev1RC6bd06b+HAZA3Ra5y62dsBd+gtkzVft/cZj7f+ZRfQd
ErZCZC2X2gE805GM8P/5WtHNMUE71yi6W3ODFHpWzSBm0COv4KZ6TPxi5L6wwMUUZCOL6NztBMSU
zaf2H4iwuID0sFVPwm3jduUJh46npJLwFLUybr/X5GAJ+tHd+NJvTpNxc6BDEPGw6eQnYAMYz6Qn
4QbVbyB8QMVM/j35fylPWQctZlo2du9koGb1Nn2ZW14psu5qUpTUCim9hwA7rjvas8xtUFKK1Bv9
9xbaMGJkzKdyQCKBipOV8xua0g3mRA37PYvapXKWsV7oSebGdErOhQyEjlml4c6GcUFhdH/WcmW+
tJflSZoL4n0mBWas3P24CDwQxwPjh720rU7pwWxzP4ZNnN13Li9U4XjWMIvH03tVw3eSA7S8zAbV
AYVktTxZkncVF1JVodDVbzG6NTWZguBpkYoY0EJ06kWKR+ypFm4CD5vlzvjAAfD6Ity4831F3sWb
OO0bu5Subb7LGuoKB9Kx7jJ9XM+WCjp232YeiQPHNFVBlNXfyR67Zm8DD6EhbHuOrxCI7rz3uOv7
zhunlJwAbwPVYSSE9y6o3WIjT+I1tobvlbpVs2vGxHXN4MKvRI0qa5D/rYBv44cUrQGZsJTJJh/S
+AhQAZ8fU4UMCk4yUAWz3KwtH3ab8fWS6294OOqPMNZ3aVUr0t0dpy4YHtZ4y4lUjM2HFaqt/i4z
Qvtm+dIT+NSSqd5Cd+TenF74n3b5iiD+vikCdgEzDzo4bMLCpimgMUPYj0WFNC1Ie8isJG8IZG26
Z5PGqs6hHHolwjeKPrzy4YflnTFNK1gOfg9dgqnWtoXTDwQjJpWsgsj3xCGs86cFj/LewnXq4DP5
3jfZ+RI1PtshzTTjbkKc7KLdFKQG7RCs+X11gwMhwI6uqgPOhcy1R6EMnqvMp7vsRxyrEy/HLGts
g3p2i+gJuER6GuAVsEBmhpn+nopQXWaApyYu2MqKyy4EiAEhVIzEI/JGgWKjTrk6+BoBwfesYvo5
1UikJ1SObTE7qgFHwZWYtPuTsguD55DT3XLSmUFOD4Gr9pYXJJTP7vs3Wp23CRfrwpONDToMlLSH
boJWkiRifIEKNl472jgBqoKLojRRcRd09vw3sleYYLW6PYazC8REXXxC37dEPNUFXyCsnPH5mdPY
B/7FaCuVIXtgQHZM6E4yJAS/wU8aom8i/GFMmd6j9wT5b5CNM7KgBx+BsMrnvb34vCs3egJLdqs+
1RbdgPDsnYNECvoCLsOtkjDD+B+f+qrP/1jcb//d9gg4s19ajJhXEIC6DNGSC9mI9POed6KRvvAU
+Ws9c4Y/lLh2E6YfnKC0ggOtoNM+HfthdA+3Y/eOm5110Fcm7dmWx51xUIUSxz2BvRG/+V68wK++
2T2OjaR19MBBamnGh0RUU1Lc6VBg8696q2Dq29+xCPhzzHmmXgKqqQcz3cNp5iafpJWs23RJ5ixy
3w7Ofkibtb8dOsIE8dme+d3VXCtEFuprawwABZYGBV8d6kLaLXEVZGnJ3qTrOT2rkb8SlyUntFs7
rTPMtDFOyIgyJtQF4qF1DhBheAUR2FMceGhzhhaTmsBXgaERkbc5OLN4gRNm5N3WNbG3YnGd5Ns4
kkJLaidDlbxVo7mImU1uQQugPMDp367fE47LZcgmzP7EPk3fyoY1XG7wH9PcYO5/tkbXsRIJwd09
v5mtOXfMt/jA44591H9012apfOtvh3kLoiVugpDJhDk5D1s6PSF7sXK5XqcMQ6NfEq/9sbYqbc8e
LkWTeKNfwLTjOOidsHANeJgL7FDr/1CeK1kvN0lls4go4InkVGnq8CY+ySR+0z+QqppH8HlRS5Mg
j4/X3GppJPxFhW86s1KJUCFbc3J0lAvxosWNLvIe9ff9OQnXfcXlvmnEwbEjJ1Rq6BWYJDfem9TD
FGVXyxoRKY3a1gsRSvqxLP27MFXbJ6Ze65qIu9lyyjpIi1XGnEsi2bcEi1RH65oX0sDXf+x+BFH1
1y6IPmA3eZF0E2LXaOgoFe6vI6PLF5h1+b4DSqskTXYwWPvBQD9WqvcFR4nZD8bGjk/yFZiNrQY/
fGS1Er4YhsKxCGP5+5YFTs7Kq03AVGtZh7eVZrutL3TeAkJvSCtJyD4+aCZGrm1ABzMIlQeqmObn
WRaOtHmmvOv1XKkdP1nUzKqq8dcU+L7+b4LxuDseNH08Kl+MXU0lTZLyXoa+sFO+qG+glc1U9Gm/
hh1TPuxKljxIhfFN0fH4BXvizDohST28TwWYwUknmzjlB0Gg88dpQK42Iv2+He0VQrKcj9aw8z87
SifNNIZequ/i7DA4iRfz6qjYMEiOwGjMQyh5DoZoMRVFSfWyvU/cTeOuK1adzR6KgPFktMLTAaAy
yHyLCIV/aQuT6ZXOFvOllKHXY0kHARnDwZJP4Ofdx7badzraRfISZ/xvtAFVnEY0RFVSqX7sONUO
Kmpod8jLTL7U3RzyvNeZIO8m17apz2iE5FbfLcUjn2nYMfDdIqOqC9dTSINqHU3qcDKTf0ZPS5P5
fEtqc8NlU4pWOEInRaNGxgjo8dA+JQyQeXDPBUr5udik58Z82UVH7v+PIoIP8DXZ7zkqLyUIoKQE
H7Vryb+SJKb2j+Z/ZnKfM97me6nlEro5Wphgq18mxFvnKsokdt62IyoH3Ba/4GwqQpxO2RJJkBDo
M6kE79CNGw8tflNkBzW/5FtufWO1+jS0YQMXTqMGduDs4uoJYsA9TU5Vt41AmdJA54U5RYaPAIdQ
Z4xhqhECEHtC15++g5dd1oN5U8y53nAsJUGhlEDD/z5zEAKRqFRQKsG9JyfA7NgRxNWb0hJXGnPp
Euu8Yv86cTxNZe1Kr5w10ApCBsqyfvU9cFDaQ7F+HKiWqyyjFda0uf+gYKe3h27s8varuyjYQudb
8QLzyKGczfc799MxGy/mrEQSMYjxZdvRAhOU+8JOBSC2Ei9WFzFh/IufBJExs6jnYMIh/+QdAo1F
Ps2SEXK1yppFO7UaPNJRQbRffv2V52l4BTVmWi+kC2r06CXG54YXeCRKrQ9McUgfAcTHQptLNNH+
Q3O+e5a+iAmPUQS+TypfZa5Jn/lj0e+Hm1Mow6UoZHoOpw1b6fb4HLl6hBPfmJM4p1C1k3sjEtpQ
Rjlt0SFEkE3uCm7dxBNMz8Qdrui8ZILJ24leF28uHFcEVgdjYDqMcLWQUmFdJzDpXYp2QICXcx3E
KN9jqPB5LvfBrvL4hY2m1/8XKTcxV/M443Lb4gMNjeJpizI4PbY05Cy7G2sljFiIldZF1snKKQ90
lw9GTDcf94W26bXUka1oRLPGx3gilsi8G1DOk9YdkyxrGj9Ek12dC978RVTyfYnEB9kL2PVn1kuq
RDeoTYosNL49Y5tkXzr4DEKGMl6H4U+22MbPjUTVlyNmbbBDg1VVgEdeRq2XDhPCnCdcmMdvXNIo
s2yZATzsYH87Wmj3cUrm6E7hTOjo0aYVRJvHfJE3JvPJZram7Z0taqreOe6KXXi/9JDCarxaZ0um
PnYwLrrA94QIJ0c4PkYsVYSAj0Z39aYinQ8ZF+b4mhn28mHy/neTj5MDUSPuvs0UHQOoc+KhOIH7
dsGSw+eQU3EARU8qUXpTVTzfnaDX+M4FPo+di0vt/1E4JxVj3G+GTTdk0ERrD/tLAJR+XET7+nCy
dJ41k9KeD4osD9ylTPqG1LzCLwHISUw3Syi/ugdrsf9AkfVf4oZO6Y6QVsfFibAHIq8GaLHggmRZ
5g9Rnpg7xoc0QQPSc9Jha63MPfZyE6yorkwK158Xk26SvfFgx9saKz8cIjnyeme9TrtOxGVFXrkw
z8UFgBtK9Mjt2w3sSN5fhRJSLZnvUPL7rte7Qe4Uc61VpaVrvd9QJj4b+q3FSjQoJ7d8/WGfcv61
jilV10T9eW8mBfENkDvaEftbGjnIsCv2t164HHMDLApthEokM8TJa/rttKLf4g/MuDmW5vKqJrYS
jGHCmCOP6lRkXdZpsGfjp4OrzkhNf1eR8msetWlNQ5jEXMDFrqURkWA/ZWP+pBwrQiVpsN+p9PqU
y9Y52rpElxLkK4iSE7W2JyeTuobVkmQ6X6Py/9BELwb6APYp5Le2l3rzE5FAtfE0VY1iq8vufJnc
H75WYxOFrFxD8ypZU923rO4PaP7MacOA3BakwGJAQq6Llu/2REL8E5uRE5bvlhZB0ODbILfmiZqF
zx7ph30daeNIAOp+5h4zJ4z5h93BlJKz246lvjmH4exaj+kIg5oI8bzEWskR2yj5iI6xNgjOlais
nhqcxrxlz6MJlCNavmAfIDjYnw+q0qCw2riCLlJrg0mvvpkmZM+4YxlbfbuhqkkWDjTKWUoO81QA
DRgoJiNkxicnt1dHYiW8FRGriz/9XGGaGzCkYEoTMk6TKygzduBWvgDjJ19SrTlkPFONwMiSdFal
loX3Z+ofL6DL0TAMuj8GFHcigi835ZYo3BIJMGJ2sMwMIFaMjx7+QuBmxc24jGLBugulV8b/MaSO
/JI1WTsXD20faoj/C4cPHp80ZZCBPlybALik4a1qLo4hVwtSqOnzPrAJzlwVLxB47koPFYbQm4HP
WcjsMzmMw7en7vyEGObLxOn0yBEngpf8rvOWCoZD9gIyBcLWm/lOnIIAD56Mi4aDSkFzJx9cu30Y
Bolh3AugjzJGA74j0NvmGibYHeQYU2itp655SFMIaWN592s/he90h+ara8kyhpbCEHB4qKtdT2ZB
cmovhPsqPJ7lrq5ge60Du9wLiwpgI/a6J2B1euDRYzFtcEMUKNcfkXkJiBiyYcBsIpLBihTU2HSm
5T3HxTJmVsDzZbQ3NTH9575+V95ROpsaEJLK/BRLEa5eCK5guc13176a7sKZdoe86k2He/kHc6GC
V7cL3INkzIG7H41bMTb96sxqF0QfblI20XPcIFxqqAhaMMK9LmU5y2qINF8uDa85LU/VimoOgcM5
h14YGQhHMRSI35DC8L5DLLunHDjh+Jy9ANB5BlIfZkL9vJ/Fnn7V07CV4p4J82rWk3+9lxBp0Ofx
UkXVriymVJNRBMiib0ksKQ/D877HUpLJznBp8X8Prk6MBjaiMkwjUqVSHCs2e2j9C7DclamYblXZ
/gRIeqwRlq0XGsI0SxgSNm0PcpDzU78I7MHEhKkQjinT78ESVvGPbBYfcZT87LmKM2gL0wKbeRS6
Qt8BbhFpCtRHwKmKAkJguHLVQeSg7GI1w9ZJ78U/8zdao9yyicEWKGeROWOMXoXAPA7ixz0r9erA
NkOjGF1HMaszgxAth0v+W2x2TKEaVTNaCAzVYeoqUOs8oO50v+fAdXH+FA+d00wAO3GSrJI99agJ
QtuH11/XoM+udBZGELy3kNvbIhehORkSQopOPoiTHtl3JK1IWKjc7oduk8HqFI5ihU9uTsm0Jb6A
J858GSpG6+SUVb1WoQWDOX8Yhcgw9UIY/n2FDuV/NAJnS1prZacKLc3ev31KvHMT4/MfFnLqo5mz
66JwqAmNeUBRqCf8D05TdOibj5BqEQ7nbWEPfVupkqa35PyIYKL0rzTXPZNGm0+Lig8+Iv1lKXyT
2yG8VvTKUJ7UvEKJiJzBmVx/jreIYZvoW0rMGHoUB5FKuHVMjR9nPF8zS5ISf3CbQb0SIQAUZPGi
ogApFplMmQvpaoTiTsDIEgpuVqywne+CzU1EfYhD7UuH3IU7rHmsnDEOL+5bdbrCBZZgSKiA64p2
vPKbJ4nmE/T1mnbMlkEQ3FcR7REWZo83fKn6l5uXdUhKfA5TZTpw+Tdcfq5bLnKPEk5RQGoYeH+z
VLjCQm+ggu6lsu5olaIHAeNcxgmHIhYeAPe+0dLUfnK2hSLfKPDWvyRf2zkZjDr36wjBFBpaHnMi
cXntaJHFONIXdEpioK3ZwaliVcUInlIOQOWZmdDHopbwzWjzAFkNPqcZ12AZmJMBW33efm+ofMzg
Bkf4+R3WXY5BsHAuWe/p5+fbhvtzwFaLXFmXy/+7rj5MoItx+IKnBhMxrdLE+qN03XC2GXSCyVjq
7zqAVR6c6ujXwZDh4kRNXNgJIw1VqRPkMnjPmCxeqOPlCfVfLJ1Do1W+KR9e04rbu5S9cfeS9889
vFVOHh+IaVi93SibFoqP779II2TP7VaSxsUSai2t10mA81oSKg1z7trRrxDz1lc9BWloEr2mOGLX
KqCMY1mUR3S3J0qCZ8hRx6kK/wBdYnR2BbMXsDFYuKi3YCdJHffpkCKWTwNj8WN8eB/hgTuzIuw5
jHRx04mnuMu+zI1pbEmqnUpyU6N8xhOTdIyWOcFQaXqphWd7+qftRyeshDJTDH7DzzdzGaCdbDjl
+fzK1+45vWZHvYf6/LIDM/lL0CZ3nE6oMWdrSARyHCyZaa+Q5E/LxOy/Ze6D3xZ7crIuphZnypwc
KBKDNuMClLiooQ6dTsGxqbSF6JoAqDA2zsXeO6fwZk5ucyAuHm+uN1E7FUqq6DEkXbMxxzdT/Xbu
c/6r/xfk4i56A+1udAyGvRpCjE8/vGmfKKbsqURhY1ZAow2r1ERHDukp9fPhGwQH2Zhw6Yw4VUeb
mi1pXdRTR4bFHeADEGPgaJkH5U4yzDZU3+qx/TZ0d0p7E5TRcyQvUrAkXkZmtxmP/bBYZwlM+FUh
Nw0YxNVQz51mNXQeAzDdwChpGjh3gFtx5b3SLAtOqEyTgi9S7D5yoWPvn7M+ULwcpEZZs3x11HS2
PP6oopTaVLMETv6S+CwQl6wkccx9pRZTpQ2ziyN6+VskTf1Q8BIrB7KG8QS/0HCplos3bEhsRNuA
sLuotLQfDSJikiYKi0bEypciayel/xAQtY2wLYSl7e7kHtccPHKP+axSg6pH35CXTGhanN3/Hgbd
HRAYGnHM+Cg2eAC8DPDqmkN/9FeOH32heIFIUsV+Eo+sHH8m7lXmnJ+48dqxJ7VuTLXCwqt8YTfJ
+gIv/Iu4XSAb7+jjnNwIKpnSpPuLPLaPuYmpW7jeDLqZR4RjhBZE6vvTKKDAss3WQqRcaQlMKKI0
lDO9ygoajYPV4T0pRyxRMEXX880W1Dkv7HylKoeTCPwuvNUEm4tIHhe8jL1R5+osA3NnRX8E+MGi
4Y9NwOO3eG7sOlrowO6ATNhAxlHxRNN+KumjtkgdMEKUpurG8UdEPWFtjKjrwLXgbQ2l+es2wycX
o6AOkMS8rLOuEk44UHorysixxkHTiUQV208EgrkwFSMcdhRhM5c4BoSCc5c7qLAtAWkdDKwFsBWp
Yg3abeNMxVur+DfsoC29o6Xv4RiWEghMUGYKjdeTFigKxmyUmGL7AcnuodShdvO4iVgDBqtXMBxB
Q5mDIungrjeRO61yuOVEZ+b4f69KzaQ2kXEYPmJ28Ft2qNn7NuBeCK4pvrWDUQKn0wnpLqPyYRMy
NTsKc0guw7gzzgtDntf1oPLbWauW1qGtoJ2frtvHyGbItbKH1XPJcOvQkTQ3HsLEi3C2APu641kv
FDC/Teh7HqNQl3Fxm5gwv6uPBJjppF1M4FEy7QueYw/PaJchG3bCQGhUTfqsMBFdI1MDBAsmsOks
1kLPLk2L3sahwLLlZtagULc8VsFJ81T4pJyqBRw4HWvlCNrpyMxpxtafapmNScmzpN54CYYm91qd
T2AtH96HKpekqWKGC9AsGdT8PWhU1MhSzwJela7ujTtqPuZ5Os+UbZf0fOx3i/GSy4GhFEAmeYKp
tJkAkaf4quCbRrzIj5NmyDiuZOqcekid1g2kWUzdiPBoiFYaFTSIFeujK/nDruegg7p3NXO3+atl
jcs0ox91h4r3XdEyHGjhu7HC4FE/iWBy562pxiI3OZ+LPf1CaAO95fplZFUE8BZMhbP70slyZgCA
1EfWseOZMVaOHY82hAP2mR0Yw/ypdBkC1q186RrUDpB4SRMEyjbp2iAnXWbc6NfhLb0EKhxiLY7G
yAAcbrEu+e3yV3IbFy7dPjSh1c4k93zKuwuRTUji9+ywyMjbbg8+SuRg/ZNgawC40lJ5CyMdNIA/
I2GUSgotjAKhfEkmor6sVKZIeAbqinJcebE0vTDxMFm32MCBIoE78aA6LBNemxtvrdQLPvUQMUjO
mwoFFcTxQ7EgL32PpnGrIxB5GRjzyFgvkzbSf4UjBH9LxRD62iiRMEiE8hVfCjc9CUvRzq+WLK8h
REXT87d+9BB8skk5ZqQoWVvN2nTVuz2TCzPXH6vihAuDhg/CWcarIGy5ceoGb6OgzdpQztxsRPJ1
vu4NjpvseotJdQbYCvj10zzmdssvDysGY+Rm5WCAff1xZFatulf+JPVhWPKJ6xq5qy4K1CwS/t9W
rd/zMJO5PGyd3UUm9KooY9V45Ucg8HrqqnCOSgEpTEdpEbfYtEI7sZe5AFdAIRKa32Mc6pxjhnMF
H9aBdyf0dMtUOqtJNnVOfjaX2gUgK1sxBl6ReugI2Hk4MbvpccuAWejirGyx5s9js6T0VTTlenHk
OZH1fo8+0xkYg1QuIydKplNmeoTpk+lg+81ytbKUrXE84zxWfG/57jQYDoVz9lqzDQ0bmdrrDNfF
UoiY5gC8TEe47OYnPQb7pP8DOyc+7MzT4q5FcWnsGBXKCEqRIcVh0yjSiZ4eDcX7R58eur1ofMp3
nNGfaGHCo8dShiKFaPlBhoHle1EHOPsD5Q3ZViFlFoG2ljFQJDYA93VtAvZ8JR2TwSETKqQplVRV
rthUMz5yPyx47k2PgZhBPuu5hnfehe3rHbNUDAjLe45qPKsGIxbCo/p7b2teFZ1utUY7GzG5kYi9
DcLWJR3zy7rT77t5+Hfaj26WAYahSbGR8NbLvvwXMVd6AZU7uYqKUt2RXZzFzoGSyQ1KQ2jjkS/F
Lm69d+zs7IRUG4YhthqiEfwICWwThiqJ1SYHzGgZ73BxU9NPWMHW44yaHEKPz5CAtbrCI9XZ7sM/
wUbHyspnB+Q72s9sBOMMiKSzJMHOAcxmNNActIgt4eVtWtRjhIVz562G+6Vfxk7KwuIl4CSpveCk
1zPJdFu9JqK93a9t0CPaAbPqXB0Mzn3OYFoemCW4evr3Zc2H6tWrCOQdmRn4YyoLj1BGHFQxG6nB
BILIOSMtiz2whcG3BDnSkHV0nEkZSpOZWTTVXM7Y7tLOAJzl2TiJEErUL1P3lK/pzWdj9c7wbQzx
F0CrdR9C3xoWSevbN8lJOqVURhkB4OcVTHs93KsHw2u4ZzYd6O8G3iBney2BNhfbwIeJZ9JhPXNa
nPoUdQaOsKIi7vpVJWGF1UnHl55RnBj4D2TKIWMXkr3teGctg/B422Vh0JyoeQV4g2pzH0hRZVqJ
Ci+VQsTr4itVlibtFswjTEVLxiKqcVVrXC5m+dMRuruSCPGeRDWpQUeSxYvhFXh8L7sYoUcIw5Xz
2OnbKjdXIGgd9oPTN+uM9ZG2y+txD6XKUIpds48t32ZzIUvsTDB2IlBYTqykY1Nh3ievrr73e13l
AUin//a0eOllGQtNoGzwVFZsYD2HBpgJxQx8J3CausiIiWFjoe5K3U9FNBXtt4eQd7/JgyXBB4Ln
7dGxGrcgm5syq88/DwYatsZAmuTSXWkty3C7poP7Ud7U/+4/cAv4qBsn+Cv7tv9JV9zZCyeKZhCW
tRer09osD0L+hDK42q/SOGvaZaJrkewYCSP307Jp2meqkNjsa6aTDvOwz1/yiq0GY1foQVDFaia+
4gCtkUNoy8smdIkASEc0qqdwpCXaEosi60vcGvo9+XC+ThhtG38HXUmzeYYbBifbiYKhwbafgv5S
g3aEfgge+SLMdPCdeyg4O9M2Lfh5xEF0LcCdi2Iqn+rujoaLQu7iXDoLKeL0Y0iVvkaYmqnoWFfL
PxG/t9ozrJGcmHrqAKgXnnoDZXxakhJrA2BcH1ayBk01lEfVTtuOlaR6Pg8RwwzHymIT8AqUYEOC
J53PUuSwWpDqIiD8aDAvrd+RyXHgkwAAymqDDXMy1Mer0VjPd9Qdo6k/xXtN1fVDFKY+/2Fhx5MG
g/UP0geuiJhG5PfL5dJheaI55tRh/gO6LzLPDm74UyPjzqsVS6Kn07NTj4J5bZP37fhoeUuwfQOg
8kUnwtIRdHNzS4XwfC7o5mi1AvtqiKn4HXV9TMrAp75+02/yMicgXH2/ZtMkG6Ur++JoaQcdx3X5
u2CRMt9dbBpKgX3K+gsWm0G/qQaeToU0cv2HcLN+MUK69XkC04/NqZM4CTgnUWNH8XyRx9cAGMlz
v+h7AYFifUNuCCTWgG4StiolpjgxWJXXeSeYfiVr1UChDCk6fMJOCRmHIZH4542xwFD1puFk3ZVF
HuiMRyqjq+EFaAcKKNj6tkSC1p5vtg9smqWmYXNNi+NK77rysowILh5JswwGcSslJnc68D8sRr7Z
41vXqA+98qR1qv8/2rbCcH+ZsBH/fTrRkwXQZVxgF8fe4zhf9BrweD3s4jUhG82CxJNWC4N18TVO
N1X8T13b41HUxmIwOm8vcSsjvx3DVd1V7Q1b4QF5m+Z+iMQ6GQb86rkcAcPA0QLP69JibC8t7Ngl
WjreyIUKeSCre9ADWQWhaV2Ft9mdfXksaWgpYqO/7HkXNWwI83u927iy52qI6RU0UeoRMiTZvxaR
mN8HDhmwJ8NaUF4KgKMy7W/ylQQkOMb26+lPyKCN+/Y/2/BS693USJDyB8obWzVTghNpzzxE18Z4
2ubB28yTg1kJXHE1lUl9T74etb2UpH7ou6WEh+MdQsRKFRnPIKfqIX5JeDCAC9pLJa17HoTTbZwX
n5R2nm3OF6dz6TAW+VFVo/qY3IU+xwPGvxn0/JL2v+sIx9I55eY5xOJDjF2rclD+wHQegXaRm/DU
B3F6bfKOt6L6DMfT6Z4hS0qGPqlGkENEVRi6KtvsW6yJbyM/6jkl/jxc32dPfI8LIho85L1LHghf
r8vcIdT+PKN+QMrroyjBhujM8UBJwV47x2flKHx1PdatO1W//5V48VdVJ+w09+Snnnnay0qpXfWh
43YFifA9LmtfXll7XDhBvgxXT/1u2Dm5Q8TiRjWQASQVFLJ/VP2Xt/Jo2j3v0pBt975HO/c9lN6F
6Hs6RlmVYrgiuPT2H0L+j07/XfrP+qwSz3kx/iu5Jf7qFtGqdo5SthyyIWdyx2hpZOsYYTstImvw
LiLWQ59tKsXNEU9k8G5Ygmi8DEkAyPzu3FGRzedHU1jnea/1oPMf4OQVNJb4kM8imtu4Z3BbQnMn
tgRB2J7+oG21M8oVYmYcseLR30DqGHmG5d68GcJ9qTGVhhtferBVCfLK7XZ7LalyFpx4vhcqcW4P
cpB+OhRA2NW3T59+JvOJ9zxhoII3bHbuy8YjgPUOY+omv2n3g1IrTD/6fSMwmshjTA0XF9w9UHdK
DNSA9Gp8WadJ/S9k4+L/utXb3BhdrOHvpk1UPMRBTdawQNUuVRYl1t76+vUQcibrucp2N6gIZV9u
XfefBn9WNPP91IAeuAuRNcB1QWOaqk/H39yaJIrcRPvfCRhNNcOruhsCxOijbI5SwN1Q0bt+emKP
wEQkgBJe20jdgyl4oO0dUfEACsN8o9vV+20wCqo6f3eOoZumTUuJPg6xJZJg1oSsueRP20QOyFm0
IJnPvAtgn21rnS0IKo4fvMuZWXOT5iIF0OKL8qrm5yCDUSFHuziUR7vaixHQ/VBlp8A03HoYu3qP
/Dn6MhEpPWJu2PuTjkoQjvhKkZMbVByuJMoyaeZ1LsymQtHct0hwJYtu8RHsl3SL+tcKp8oiVq4q
jbNgOWmvwu2b/c1ST2x5FYy/Ml9OT+FNP0r9L9Ax7DknIRwDjNETVQIBCzvC6Ye5pimfmpGY3Zlg
sWpceFIEM1IROi9Dva8n9RengORJrjL385ltREVYm22ZZ7BwNLNaqxH35bJ0Lr0pleqItfIUs1s1
Jw2wnaCFHIdweBQpqqyidhiACYQsiKRniiVkE4b74UDhzfljqFlzCdaHjFySYlWDmS8GqNJV++i6
8oZUH5Fp5XLxIf/JdGZAJ0+8TtdXcInyZGOjBAh5kxwAq5BaI+3srAMzY8lm1z1kQBhXOrIQ95T2
4lgxSWMV1Jy+qXyeWTjnrw9xo7AD9oLL1hT6eQehhXhjITamoxhX6ah4Y4S4zGJvsPaXNeK1M6dm
8SqEqtge2e3Yx2fI0NYrmHgNZddY1ILHHevAq/7B89wTs/NKrTIfnufxD80JvJB+6JNRqqiy0RU7
1nlYaMB2Ui9dA70L6JwdokanBwv/VqaMJ7kYobQwfo8LuCfMbHvavf6bGnRJx+fl7uzUQtVjE+hQ
PZq4FRmO4EafjFqAiM66YsMR4A9AOwgS1Zi8lv6w9B9fOf6YoVuOPTssQ9baS+2X6dFu6j22Gc6A
o2T4St2UbawwCKsdrauDKIUDvmiRR1zoB2gXyn2dnfROvNMYQs42TixC0j4uv5hjI8KIGAEv5xkh
UqvYm4Ux9sYIhMG9CnCH5l61XDnpB2JO7druoiKyo/MI/4P3dzNknGFH8XDupXIcXrlLqv7lWurp
FhjwXM+w6o5ug2hdz/w9Ex0+NsrIDaNzLXkajAmEDfqtdMaLZXfZ6vwQkKEzFfbeCC0h0hVZcUrX
vteogT4cY8EiMoyA2ocYrK7jNJe6OKQUGsJQzn/YcKvhzdOjhHzlu0xIazIfbqlxNNowmsUkaZvG
HjqhKjKq5YefBzLxTESMuPzBP3SpS3TH1zyZvYU3njwxlnTmPRD05+F/jQf+T1WLBmmXlyI3mf1v
7WkyoUCyb6Oim+AIwMDwoDqS7lHtENOpwXAvzsvx6saV9dWQnARGhtqZSiFFfv/5Ezxc4wQOCCDf
aq6Oxy+6oqpyHvNYwPX4KcMM8zP+cxfw0Gtnru9B2zZwDbzkNh70Nhy+AceokzL2FKdSv6qxjOX3
X24z+mMtmdEy/HK0HHwAkBBQKhozV2cI/r+ABJyS2Jt0yh6oO2300WIYAI8y/ZWYq6ZwPOSDj2RC
qj3hZO00VUCxj524pBIDCfMYazNtaKw4c/77IQeU06g/GARk/r1vQKG3edRSISLjBj165ptP/TDw
YAZH0gGprCEbzxGS8/8m1E/38vIKQ6fLzPQjctd3Kjzozz46cvD7K55hjecpTR7DDGfSxRleeWnY
DUXsb0xgkmSbK3t8sJ9cQ7n06pAzgSBcKgWLcaGG4YrqaKoY8SMDUv5qtK3vrF3cgAcuWb4lGJxl
ZGpaqhQReGUoY59+4ZfHYk2zcPYiRpbfuchObQHATvf438QfIeTjuMVh4QXFlXC4Jmch2N06Fa7m
ruLCo3L9uV1tDqfW1WFpfqRUGJg1z+gRLPO4T0S7LsEQt+6Rg9Jbbz1g747y4Z77Pw51QJ+5y9/N
1K1fGU+qBRpZNexvAEWiE/Abg0FnSK/mx1fAVqRcAdNpNNVYsrPssUxGZceXWKhQiYsSaoxnrPG5
/vQgxTodTonlJFm2ZYzyAwbRADHpdVveXo/TEmLSyKkxzcD6SDgx8B1dVC+cOi2syT8EvmMAGGbx
jtHlJWnljDHoH6vNEyHcIYiKZzBHWPhvu1uLEcZbSarGhR3iaif1fCE9Q1Zbm/GZJrCz3ASSsKRq
a+kReWUIgYgdwyuX17yVWJSukLQS7roSpCKhulVJY0eYKYwR77jnB7C/uCYWd0elA1e2T25Infsp
VVfDLMbirFPZW9DHUMbAeLLA4qai55vMlgKGW53OagVrjJF5SiKqypO33WmBNzy4TCm9j7vpZ3CG
93H10Uyhk16Po7D5CXkbnFzZAbDL6K5kW5/JMw38rfpkmNJgiKGFA7jJm5cKIKClDpUrpLPKQTue
zWDiB9D3sVjf96QdzvdQeBkcRE9+xvgnpgfansHjb4E8QC0zDXXMPRNzXEtt1ZIaF+tSeLBOVJLB
39nql0EqtIN6VZOms2NyU/yGtlvvBbgEHWrLUA99GYHZtRMt8/XfvGwOrrAJ77cC0da0FfaAra+J
pbF29iQARlhZA2Abnt1vrR7onELYfd8TLNXix1qGP9p4suLQB+Pu+guzVKCAg3BRAUy3FyYtBsXN
B9a4BwE1W9W62JXsVk71QgN354VbgjgepBTntbPA7+gKD6w0/0z22VK28u94G/E7zRu3CVvx87Zi
LK2C1ZloeKaVU5bvEB4U+PkOY+AvcPS1TLjhKzBO1D/uF5ZjV9KcMxq3VjOHhXyVDmWtsziVmbCP
mQmBiWB8rtJOOlipsnxtzFNQQMFfxJdWh9Vz9Hk/gO6ap8M8gFEqzOD2hBrqYotKTi89V0mDiQ0w
ljjGbBif2H4biPR9EDz83X8gNKPJmqYFUuKtyTWgxUCSzlP+NhFU7/Jf/dzEQk1PhPa3EnRy/eFm
i4n2EYLFzbr+fozPKw29JtBdav+HPhr7oQTAG94JEU0ndDx9ZHNV8AxVXJ7ABN2XpKMOyYi04o6K
DyXQe3Qd1mjdTxOcd1hTpdwNxW9fGy1lFAIPEe3r+a9M/1eNSotG9e/uELqN/cr8vvNmRffkuzpg
DVgLEx1WWo0au4c6jP5AcPhj8dWRba2+vH1VQ1qR4no4RoD1uchZhjtZM3SaKzzU+LsCUy2MEI8p
5a5UzQywY4wCvsg7n7fzxTs9Xuslgm6VMq8lXfyvHND6CcNz+2cz47yyl+e/3e7gs6vhBaeb24t6
7SogJFcSiS4eET3aTKNn8GPfbg7EhX6nXes9GESbQujhtRyoIpeNtZKWQVQiePiPe2DLJ8DkNUEz
CZ25ys1KRUnFJIdwXUGshTTvWD29O+agw0ooiH38EML0BmJ4fuDT93FoaimaPrEDKdV66hYAIx0b
WwAbuQ3dKjgAChrf9nNEFt5JFHz//fcLxLwGDOvdYU/fYABlS7F5ZaINNirl02vd00l/1b2Mql82
Iju0MD5XfVN9yfSDbr+zUNlkNs4pku8gKex7NQLUELqki/4uKSn96JG0WyVuPzo1273xlK+GGwEG
lvMTpvSQRJwLuA6rCUQexpNQWUmPI6AcZyph+dipBMFWZBIy0yszxaiLfv7ziP8XxfZ47v3u9+C0
bvEpH96Whqek3mxOQPZudCJUi42o9p+dS3O123o/kXW3eh3MEbZFF1kgVCkz6uouyrwDytMx/dC7
ze/9rqKJ/fm4YG0YgBurAmHXwpR9Kj3dcWziha0/zF/nnxHsjJTlphNeKXEjunBotsHeaO4g/ag5
9GukB0gl6frMtSgir+8GANoIJZ47wt6OIlvUSuaGE3b4/Mc/6piJ1Vbk1zluAWHcwTguBC9wUwGu
R9JC72OZt1B+WicHCrGVa0CP93rmFwhtjvbfVQkl5+hJmP+o6mFn5VqirBcThWl2INqZJ+99xk5e
0Qi2kFkogvb3VfZzUBKOrBymQE3TvCIiErSPUOx4jq+qfvf9SATZT8EJBtgg2fCuxUPsAFjbFrVV
znGt9m9zcG7TzoodRfP/zr/zQzu5IKI8t6UmtdP2I74t8yQgHxCLxeni0f9Fib1lwMatG6ftJ9Eu
gDDVa3PenRUJnZ7jNyk9XG8L9CyuUWVXFyx5fgdgHUVZfO6wZdJUkSKyrNcEfbAtY/g23P7qgiTy
ShTvU9kFgEJkgbbGA2LtMQdTuG8+wGTPa9mMnvsFIl+XRdKNFwc/R3isaH42cDvlkdPwRx3TjLyN
lk53V1+/6drnziiBai6HpTNAhwU2q+RJ+0u8kNLvOEWwzl6JQCyb9ldMaOMKY3vPlXZUWKhlOmYn
DawniTCdG4+0iycOLVuLplLRDzkPeyQVt5k0iHyUjd35f1wRvcl7uq0LUobWeaixIddyh/85JDVo
iwjtRpqUPH0/M3Ngr7wU95tZrqaeA86i3Jf4ME5L0kSwSyqTUsROqeHUkC+ANoJdH4Ce6BnKG9iO
0q58Kbj3RMtEBb3itMJyuoZ0seh1M8xEsEw5HVzdOsFnEvPmNiUtHEuMeYg5y/rGRQhyw7FV/Saj
eznyyxYJFah+iQJAuQFLel+xWDalw1cyVTj3aHP2PYyF1DHwAZeMxpPpanKDepmsVGlo/RIkWbRO
dR4eWpjyEas+MDcuhobjrJ537dVmH2s7j/qBLcmwiI0RKe4ljgqCdNVPs9aWn2d6Q2dMZ/0Eb9MR
KgAI+T7FxEMPzK18T2pFJ73XQTEX1pNSI78Wc50n7dbdGUzqG8ZtytmtX25HuqTMZXCzoIuE9s99
38COh5D/nNcjNKTH4IKDp6UwGDf+VMYHylWpuyIiLBiSB8q96JaDy4XYTW+3uW/XY7yB9AnlZwQa
3Iv3zmB+L3HH5qpNiEA4uDkt+RSiqJHQXEsbMjy9/XyuzyMLuYerKDMrgOOu9o1dWyEfvBsX+9IW
tJeCh8teY1B9UN7jJX6cFkfyLZkFbJs2UIXlQkoDSNTM0fwcuNVWQulmKxEPZ7sbQaDXDc5kdpec
Bw6LfqMU2Cd1vGvOyqj11cqsWVRuPhwbRXtWIFZM4vSFrygB2epMofFPTkbzqGo2U5xma08dYF5c
VMxFFYsA7jt5HAKiLFGGeDD/Icw5QtpfTRYCYiXrMYI6FUraM6bpe7RcRAkLdRQ4JH2gy6BbTKpU
tZT6m6QsjoMHBHSv40pjakbS153kPXiHkJ4mGcX1MyvEMpbWHqdeE8FFN8g+TVn3EF3pd7JGmmz5
eQ24UYn9ziyNd8YiCP4qvAy8iIrKm7AHx79vRRqYv3CFQAo4wwecDiPSYSdilTfGvDAEteMx++6U
LMLc1Y0DR4KWvU9UJtnBF7cvQUNo3ylOa1cgyx8hRzcwo3gT1DFhMWQzdItYAmlrxpD+3loioxHk
xXb3XTP0hclU2BGUwoSe/TrCyzJKpzR5t3uOLyzOPT93mTo6NdFtqm2EeD/gfj35IeaBYd1KVjI/
jlwac/xoNi158xCjIypu2il+W0TVySK6DwAezjAJ3KdT0YG/l7sQhmtFJhL4UUn0Qqr9Brb+f/01
bOM8CgZ7jqLjNWurhuplSQz3DZ0Z5awd39Ea7hGKlkzG5m2HZUYlmftWlmHLIBpNB8YAryT0iBtl
yuaBk6IrRIxOp9mU+GCkWO1k61iOrlUWh9mnV39blBXvFRuu7RMV6lBs1MXcDdb2qX+OSKOC1Gr4
lkEWUbb/7GlogLCTqOdsJwOAO5FBPMOHqApJZSHcsEtJ/4hOXWqPVSTfFBCsNMeMK1XDOQTIEtff
vxnoQJMzp/eYXSIVEfKp+/xfoeXZDiTYhq+03e3Vpm2XJUrlR9s6vmaFfcZW8UYRDUwN9pF9uj+f
p0LLKrMYOWPwe+PDpMLfbjFY9PI1/H0cIlfe+oyqO0KBhhBFU7HoFsL3155TNTA9VCjItpzmUNO5
i9HLuIxc21dvEVQ8kXberkxh/eVaFdcVLmFYD6CKCYkM6Rne66s3TOlQvs+O26rn5okd0F8Rx+tO
IzX9Xxdx9i6mMNsxZM0gsHuoGbpauMbeHH2i8MMxX0xuJSmPmDIZAj3rGbL2v1XaN5yLCZa0bFYt
ZhvQE3IhnmedNcB2zcd+IJB55S5RlzSOPsbRgCfCvKzsveQRRb5juM8Cij1rAGWJt57XQMjF2fJh
ZdvSjZmHu6GI8Jc5Tm9w3MgE9GQu6p4Pa19NuBJYy7vak7GoPu+t5tjvXv0QCt2de0xuISTXcn5G
F7sVVJIbOwUdxkBaJEYvZsfBqUttQhsNpEd1e5vuL2cPBa2llNEyvHBKyI2+EyQjLx92Qr3wS7gU
RxOeVh1FYuVCGeJ05D6VH9jd87/TAptrciFJiyYkBjWDROG8ChoEmXa6Pa3CnqCU/hUNQswicQxU
kKJqHOOmFoHjHb4aS5CRqJuxCvV+BCKjyzm0AyEuZOu6nvxpmdpLdk10LudRlnoSkf3fPNN01G4c
xm+u6GhKDnxYw+/pCbLfASvFprOpYC1lswTR0qMcFlGakhtfMFutckBvQ5Rk2HNF4op0cQuurz3P
Vve4MLre8szt+OYS/PhKcTWh9R5flWD37Z6UgksuZy/Fyw5G53R5korB9h9F3ThXSYGoyvTa6P49
fZ3ihAi4kTmpHFSii3ngwcOPg+MHYkzpCcwDT8TTcW4iSKvbmgDRZSRvJKCaaVvdyT/czckEuqw1
dA59skYQCy6kastgavRP9MP0+2OkAgWjkFMFNfmdcT0alc17CJFHpFUGfJqhGK3+LSxRnK1zxCUs
C41yJ2NHPEozbxihQxJrO37DS4t3SQw/eQabmipkMZhCQ70hRCgpJDZeN0qGqG5x3LzQF/tzCCs6
7V3loW23lfV8s06mUVCPy8hltVtKZqaj3hVJ3LasG2kQh+DpSU7maOvwwimZyKXz+dWnWUw9ZbaM
7n/QKXWdJG4I2o6wkIc38YRg5GyxNA0SR8GI6U4AuXROT1jkY9qh44vBJIt0hXp84sjf38XLZdv5
TNIPGu3FvUR1BQLNBNRj5cxC8JyagodtwFnyIEwIbxFU6ewcaMIUt99eRkZP2IoCO1/tugjFqtxk
8vWmztP3KJFf8NAH4+XrkxW6+ooe1MmKmEBjJQsD0NyPmhCnc0jmUbBiX2N1NlO83gBL1V6t+J5z
J+1tkPUFt6U7i9Uq6N8s36jhXRza7e0i2I85cEJMldvEiPq0d9TkFDJ7PwRbCgx868ThwbhITqDx
iDhERnp/8AQ74bt5LFxkEkhwmIHgYZgUCRVZBCIMDd4Faj3P4glpP+6ML0bK1rXs80z1mfUaaxk7
8cdLjITGs2nAxzaKucOfJ/esmD0Ss9rl2oeRlvTvmGcLJGDel/uzOOkOpfJn7bmMpEKO5rNl62S5
cDDwyzv9XzslVW29ool4Kbso6f9SsY/lfODWiZhAcWMtoYh894/zKsLtzzIho9/Blr8j7kRVStnN
AtRhxxz0/O7YduWKlitMj/6ZZXeVkYJYwYn1bpNhF4JP8yNa/LoKcVvjZjxGf9WCYyl2gIznIX41
3oFfVgk91/sazQTOzvblJUMEghkdcMYvOJi5uW8ZBcETNooHTa2dNHox5fh3UOyjnqY6hGTKaUAb
zhsAELuFkaCk2yY7HiXry0gJDEkbjWi+dXqgnig+OAENljg4CdcScDRzJMfS0Nbed0pUS5nkMYym
aDcJ8VbKTnfc9fu8Mw2IsXE4aLj9XIZTFF71fqqHJbact4HuKAr/CqwO+T9bYwUsCJHDDBsO/enr
7DLQkh0ZnIm4TGuiNHGw40dESJt5C5RSvZdG8l+T7XCGWGcWy6ko9kLh2hidzSCJk3ojMBv7juuC
mWlHEDfJAfXkfL/H+SwIry/oFJS1tU77CPbmTqaOQMNyEqGt6M9jUsOuJPlvudZoFrNjBgyNWZ+C
E6BbD1Nm14X6y668PY2wveVtwDIs7CXmFgvBC6I6V7ku5+Y+CUgyXvSye6D8qfYpyjY6V1qbR+JT
fifkIeadyeHtL9Y7UbYbmXN5eGFCvvYwXjE2LcAdkbqQ50fSIdNQ1s1b5hgzYxhg2966IxPG38P4
uUdkUBIixrEtTNPhnpYU5bO+0XF9g2fTA935+OQDMlrEgEadanM2G3M/tzuNhK17HSCT4Of3d+F8
hdUrwDujZAGtsLRW67kC+kiYOKJCgarTbV75ezVq7gpQdZvE3Pwp+j1Xd84wkpztlp9tjhbV8ULm
u7bTR3g6Lnt6rTwvMjmcA0g7SaP3qk4ZI8WqhQKH3zn2o8yb6oSHlLF8JtcwHjw2hW199zH1HAkM
WfQsUHv05/jO3BC5loapHlzzmM7BW/s7H3BZZmP0x4mLAxoKtryrAyJTQCuR3Y8Hi/mbTpWqnvbw
K4HY/vdQiTUi1rAVvVLQrVFw01eaHGWC0fgl8z2RGlMpFuRT4AkdgEYYIlzCCMemlQ8ZV226mpLD
V/yK7Now/hB3Uo5SBNr8ilshuubmOuuelM28zkXogbLyGQvjuhlwuKnxSfMc/hceW4gSEF3b5yy9
R+YCU4YwUWKV8g1pnbdpfXjMR6Agd1fo5Kl/8MWimoh4lDJp8w5D/8DzwLNqO0vzN7C7KKvc+Utg
lL2JixgX0EtSxJF03zFMVsxvdGVVvReZdu5QVgPYDs+/H54fQECxkw5FinNAs8dVsPkTNKjFNl/K
aZ5OjILAP0V6RQG7Q1YdDZ5aExqhNB5A6s1L/m3oxgef9tdA9q+VUBCZaMWG2GtM+CZVXQG2Wc+5
RfQf3G7JL8urBcJ7z1g656mtY0xU4nxe0zj0+kpyeTUInx59EJFPqu4nGLAz1aBGeNT3Or6arrWQ
mxt1ijoQEc5F5pB/uWH/wpR/H79fXyoMHwvDHJvSwxHs15+pJ4DKmKU/YIQZp6g5xTzSArfS0Lwf
VRvJkb98RE0LaU4PYr3tRrhNKOWKBibGsZ06SYF8IjGi5qdeCL90eR3EmpGmu/YUybbKmhWaK6iX
SdmQGeF4UiRUHq8Z0NO+mglF31xPCLgtIx1bb8BS+fFZTA0RB/Ze1vK0Qn7wSBTuiTq8HODPBiSF
pxpIYy1ghYk95jpFF3MZ0XNqOmnaxp1+p1jvpowBAiVugXDv+0FSargwX/UC64mQd0A997qqzzfq
WTbZ8WnrQj2hlHGosrkNSnj1bTGJky7NURRLDQYEHzmhwbLUeF/CqYpvNAyrBkjHnp7snKlnhEib
g8vXvnzYc6fC9CfIrlvusrn2vG89yFg29MJ/JGN5kg6ftA5JPDI1OZGzELZYQqkqiFQdde8kFN14
MxMUtfMFic5uY4Pn+yKTEUpPe1FhUZzsRAJbyVkh0PVG/O3eQkcmjHFVcH56r/6V0ykcCN4cX/5x
J6gmAWKpSCabfvbfGq7NAC0KLZZx7aEDOaw366YtnGFWhvVeIYacN0Ke1JbYMvLtm9l0/9OqAcAD
3MlCVCBy2QIEEvYT7ZCV4AYnBIdRiNdBwJX2zK6BsV03cadX6+qkzbupH6V519G8Lefo5lD1aHdH
r+ZESay8lXjZjzMHiGpXLmCN/IX4aQeQ1JpuSnyls3HS16ke0x/+q28E9dDvkDkvDe8seZelxxAv
4WGusaqxP+zrm/IPsTi4poxERChJRD2LFnNvSMREp6Juakl4N86bHFQbQj5z1GSvAZEF1CK/9jV+
VpHTHR1QndLL8poKxrEhh2fcSIAUjJCvmqaZ8Ikv67JbwMJal0P7++166fXZU4RrUkiXaduboMDP
WFmJ+LpHOhmCg6MiISS7mfIPwosxiWLWKA9kU529jZdT99cxMjUp7JNE2Rck6z4KrybCBaJTx4bt
PbEIWZdJg3q775XY1UL1OsVb0jjOLwYkIRLlRUsUZEq5/k5ymxnaiSOyWGjDMpN90iIq4LsCZoyG
CADdCiYRwxHdId9MMGnK2EkOUO/PeG5gEoUCtKK+7bJdpKHnXDbMQpiqLv4sz+HCkF34p/uJslOY
g7AMuccF8JDIUchCHA+SMZVJrIMFtg0hVAiGkIGfVW/oxd4Ucx+De4gkNQE1kZsZJuAoR8diIdD2
zBj4lKei4Siz0BuVFMryh/zj4Owew2tMebBnNXO7o2jS2WVkXUgLubKeeEwsRWo0pUGpovW/ksa+
5gKoUECQE7+oBLc2HXp50M41SxrfAQnRmu/WQNX6MxhK6r2DhGTTBcqDxOQlZfnADG9/oZ+NY9N0
xOh8OjtPOOh681y+eOXSjLEXDcafdVAvfT6TUuFg1brSRWgzuyI5ZWuU4z2P0U8L0JsTzAfulICy
g1C+Hm/Io5QN2dQLJ9G+zyPlo05jk6BMrqlAwMRXSzOHw+tciOuWH7RoWhF8bA/GofNKtDQl7ASU
AJzTm0fk6iCyGpXwpTvFM/7E6a2V0xH2Y9t0J7y7c+OfjzkyJd65VJ7qZThNwbuVAKGCgPgy2vSM
y+8/gpS0MQKqinrzeTZtIyBBRIkM6oKWh7XXq5oC6nsiJwdtsGsZ/OYx7ygY/H6++A6PyHR14CXw
PHfPMpVm9e5IG6Czgy4PX8mYqPccOr9i9D6OAyJn8R8T2GV9r03tKObdjFSRqUXucK78lHzL2p8k
/E7vbhWVjvVjyRIMt8D1MWj5zdp0fxV9mRcDE0Lhd71ljjZXfAUuc7I3azpc5+z2GXhF70LNjN48
4WbY+m54WtEYFJBaF8kTRokUiBixT1tAA9OgUus2MntzfQRODWQ2wKQ/TVhUTFs/jLmrAqaejkSa
x/Dlu8hse0M+Vv9yvg4SKRqbPDPgpYmvcbsjwakv3G0MwMWify3VwQt/iIw36i1f8UqS7/KQNTCT
FxKHp5MEJAsvQqjd7y08PTgpuEY7B1LPe6o9vGUQ7329+/OCdxdXZNzc7X0u+lE7yvXrYan61eVt
e1jd13qMtHjuTEhn5586Fkda0nsFZfwVybfyokC3oJIVMwuzxLUg6QXr86yR8NZqv81umSsuWots
lWy1BSg2jrBWEw7ZlekhQpA/gJQ94yYk/b2nKudWlYiQwMzcshEHlYCoolksfNhTi2bohASAiLW5
t29IpcqjH4cVhaUsnRZiozdiKp8eP6QHbYfZY14nIXccw8oMjlqiVUSZLUCeNf0eBy8sDiq+TRZd
RGTDBTGGK2lo/zK3wbk9MFVeST/iwxIVgVRQyHbyIALUOo/uBKrVvINBjwOmfWksXkplIJIlQ49W
VtyttM3o6U6WXscoSUrE9BnUo3Mb9563RsCmB4OWb9dlmALYjmH7vBRBBuxP0g7bsoCZ+P1N+PbQ
KYqw+lEB/iIdOsDYJYIGQoTPSumZ6yS0cE+fN188fxytsoQdX6KGJno+VSB/10tjdcwiBiIJC0U+
caPNw0uLodL63VGlhzjdD9/IlBdqenigc10hw4uD7RChW9d90fvOzZLLQ0I2ypmcvKhsFE2+O+j3
cDMlYZf07TjsSr3SvSnVt+bYwRVNRWaPO9LwzlVGp4aOULp+cxFVZfK3BTwQRmRKKT3njuGJoQCt
Yh9ZpcuYxhR9B4rzn7LWoh6eLRIiPyPinDSbeBT9DpM0IyHx74Z+BBG+Ekc3xxfH4dQ8ndrY4i9/
exRiQrevOua9NzNWOl3PQ7S3bRnI0iU9bCUB8N7sYGmcUK4R2h2nMvIsVpi9vfk683JlHr/hKUA7
X1kRZGI57ibV5x4EQqED0cpmTZCG/QhXyU01/UkSfi8DdHpkz0NFOhe/kBWxVDkGC1r59uTBX9x3
et6j6VSCXShqEnxh70Imxek+0nZ/BEeUScZY79u3theAMCzKafOqjdnvuwoxIAh2UCYmUg0BnTN9
nYaKI4MDkY2nndhKQQVZ0NlIjrhk2QoLFxWzWyPdzibTce9TQfxohHj6LhvDGjORYsMZfTB9QIIk
sL5WabhqX3Q4IT2Z/X12KnFIRAm3f38n4BXKxODcSAdLhOZpOhHoKCrRwekFDcksWubHwaQuypat
Q7jLLaCztuPjIOfPnC5MWT2vNRLfXLZKjZnQU5I2YhXRIlSZtJjj2rWlsBEZT3ZeJMN601Cp1tz6
3e3n4SN5c0wt7+jEJKmtwogPjJGePi7EvdFEjopWEXHZ65nRY3I9fuTODnauV2rW6Rsn77aDvGU7
tShaYdgErihHdzwTagVrI5RO0aRN317pgLoN4LUaVwGgQBomQ5gM0RKnKvFQNWaOP2DqQ8TWDTeN
vYSy0GwxtMpTCYHTjfDxCeQYo7JjCp6qS7WUv9JvaGu3egyUZUn/DiqEq1VlXGdNavg5rmapaIxC
0JzUQMUgvacHqnIkfG9L1Nf8fu0lFsGJYZD7vktc4Fmv+PPOR51WOveJ32kLcxsrDktHIG2WBNnT
4UmpkGLTH3cLUSYpUCFJ/UOJa6sM9AQbgJGvjYTBJujx3VbxJc9UyRikbbrXctLIKJrbwV1lkxqJ
UdZoJ1NpgLf5DA0NZPsmfdee4+/bGpVP9UDX4xbZ8qqoJWADl8Svhf7iedHxb8cIo372+bY0KiFl
IUl3OyIg0XGS0Po/PUuUy7e4CXYY3IajiD1jBoyub1R7v1LC91FNxXux2NSlL4MU08dRQP9BsO90
RTxmhONoLSPZZsI/CnDjDXDIOSfXmdUFDqrWI4hXgExa1sQTji+2IeqgTmYfp/NOb2RPDIv3asNP
13t1GeudrtqdpK29bI8sr6ycSIlPaXZxD5o3HMMHiOXrQyqaV8hTf/J4mpssMJnt9lBd8NbL/fbd
n5VV6wKhh4FNKhsexfRDW68dWwr4YDcHyidvuYnqC4NSXhgVSFFvsGKSYbXY9ePBBszrt8yCGI1y
WO7tsdM5EKnf/E4LWqDbcHsmHdruFarVIUMQlplXmTbLjlrn0qQWy/4N+jR650ny+CAjaokVpsxK
4YyQp9w5IwFtLnlgdt3fiq1bOUvq/0TqFlRuWIhs7kqm3JIes1d8IyCGnZ1IHof4FF+AoUyxp/UB
a7hRC6mr98OH7krpIbEMZdCxxsmW+EXrVSte1ItMLVLNuZQOJXij2kW7B/SLy4JfxfFwHOm73ow6
xXSE10nMfK6/jTd4mB95WEzwOnZxIDjwTVjJorI0J/RUAcwGyyQNh65TVJzGPekUKE/LFpmsxrSM
YiRdZCD7KLoElFz+vCrZzjwva2kVRV24qu4boGdXSvtsXD23Z6YC6xZrfdcuq/TDZetGPl7eas8l
87Dj2b2h7HMjoOn9+5k8B7m059mQs3ogPi1uZkG8k//UlKl80vJqYrXurEk+PUUwMXb5Ft81vcAV
gtc/PeHjqJdtO2+njrBhP5PW6P5VAPga2sd0nHLQfAQ2DDzSW1l2aLU3XeJzlqSXzEY4N3zvL3U5
UhI1NUsZBzCK2IG29lxnOpsqmCSVz2jbN5ekXv0OxkFi40Bol6M60kQ6BOUKM7P/hQUOydvqQiL/
kLWwkrTnfzz5zIpTunE4nw5zvvtYiM+j2WBOGP5VP7QsUpUd14VDhdcDKK0mY5jtHA/qRCHr28QZ
YA8LrNlT2aFTvVGEemvWs6GhEU99aYzq3LR8c6zyWdg911RUkFXVVh7t/knfH7PvGwhfPEbBAJVP
7KaZlA+e4mYmWb1JLefFWFpfqHShrYxEKo9NkvLwsJKdbxkMUOEGNKpFcAgr09VFXuNDCGXLvUce
cImcGGuR59v8I6qn9fR48SFomby0Bviplk+rFMOB3+3ZGV8nWpzHURwyiPVpVVdaSghACLkoQ164
RuzFP223MPzz9dQlqKJbGf8oIOdE5OtotBCyKnDeEoBj4n5S9Y3vD2TcXt0To5EwwuPJsNJ2Cmn3
W3J6zMxzVL0EsAOvAW8YdBp/D9TaMW7VQtP29oqkY6cgKFwdw3rlIu6qGF3QeYJI7Lu2twsKbBh7
53AmiccGaoA7N4O8mbyQ5H8ne3Mm4dvftIOLatf5/7s//fSRclvJiSvaONQCw4vnigz/lIEk3Vdh
3pT8+Kn+oS3W6qPomZyCtnyV/hPE2PcwwUBOXk9fBpzGEFdk2QJwoxYQ2geKDyfjJRqZFgZV3bKE
QBHaLEn589Zinh7p5mUOcBeAZDr5IujL/4sC9VTbqUVu9hWHIyrTvOecsHQaW4HDTz9FOJlMwHGn
V2NTlD1K6G5BQSp5D90lebNRtFO3qJgtmMk7ijpTPJAH6YQwmPrw7CdVrSGTMfE032tSDPu9Gtsp
UuMjRMwcYU8OX0gicb+wGCGfXeXnJK5njHFj2GmKUSqXss7vZR5bBQMcWFK4a5WStKIuNeIpzLnJ
3HuM1qszrZx/FwJ2slBJ5RF3Y2mQ+0K1xeE3T7fDiUXFKu1snjQ4MM19JXznYzEdKARoAL5qlYco
BXqlbx01Uk5KnSajMp/tSMdZ64mDT8NdrUTK8fTLqhIUNbBSFnAIMQhMsBcMr/3vQ3mpWFFVolvW
MVNOaa2kLwc+vuCSdhTJ2UeJWGLY8OafXdbP6r1EJ2c+uMRUs/Udw+kY3XS9DOCphPNzQob3qi9r
PrlsKi9UEsSep3uaGsa2ek+exrnByWEQ5/Io2u4LqJsUIHd9H4W7oxnQo6lzWYkeAOrYJNxx0svO
TRRWvxlmEv2kH611ipiIfNkoC0mkV1DJiazIbwNfeCFRc6Q+vBkJsbjiHjsBkKGnV/5GUn2Sfgiv
QSg95qqMiAoVmdzUpcfa8Fe69nGbRF1zacqU17I6kKnYLNVPh55ic98dWIsQN1Ld8bX7dPurqYRi
o2YHdiqDC/hK+TJHWm023g28PMZzBpmb6IyoH/XO3dv9QQ7eDswFRc3EnHNm+6gVe9ajBY87qzv8
19DsBuLECJwyDqOId8ay9TumEtPw6+fSKU3A6kFJo1Ky7+1XSVcUmkVOVBxfWb91UfukeTO9MLKB
1JShLb/6Ow61v+vkcji+A6F61pbwC1SwfrvO6OX+lWLRjxS+gAXJVrZShBuNRwsyU78YHkXj4l50
vtu73IJAFFgydB3ZXwQGXMnZOQt+IrkXLH+dexnjq50H3cKEj117SCyV4motC+wReFZYVOmXnZQB
rG8hc/F5/R4+p/qMH8sQ6C5EX9HqadVZqUd1LGoBXW3RWRLGIDlluu7b9Yohp5vM8uA5u+ddkOIP
RE4u7ODRAjraq6oUUopQkn1Z1R3XpxuSa77ADyssJ7FlZHBBKD5kSeNOpad01eHviU8qSq+nXiXE
+A4wDgj4rjGOAl3fPrahqrnKHO0zLY00ClqeKag/awkS/HGxzJ12Ab/JN+fmhyhtPAvuSq33ItQC
phAy4QCscYPBhXU9yzndtSwuqXgiieRRlYVgyGU0dab9RGsiOVyx5KabkXEljnoBvzov9YzkgDHe
NGRw3lDozMPZZjlgJWeeKPmZdFKKtnXyW7GIETpuIvNy4FEzD7SMjN310jJwPl1Xw8bthVm2ojxQ
wT0xEMArdLiBm0GRg24CUpQw7BMrpOO7aMNXuM50GlFbpDUj7Mm67Zi19JB0ZSdPiLChSlQEdQ34
A8J9Gx88gNGPFEcsnfeWnPwwrFwMUXZkG5c6k058GKs0oOKjkGXO2/xntVabp9Jpr98C8IwimkDw
pXxPss3aEBsUjW+7Pff01TXkJE/3sKvT40fZlaBA/ZAVu8LSC+0NJydQUeB3VkiwVxD06K+vxQCG
g02g5Fg1KZtVGXYU0Ss9zXhP+E12DPZ7rWw2nccMHU38sR6PBEXK6SkZGU2ugmPc1bf4bLokTYoP
iuZ6nwEbJbEv/0AAxQ7aOT3qkHebCDWw4G0vyWdEKYixc11oB4cpaml3LMMyjhmvoSOkuNwO9lSx
9fdxeKzXrfpsnjSshkezrDYhIRy8Kv9a5Gq3q5lpMrJHx+uNfIqccmo/DCXE2gbhCoI69hlt9nPx
CS7vgZyPfF/u1yTOr+CgjbovzeKap+YL06tdbSAsoymGOl2YF0XlEMyXYqsg3PSOn5Wy1fa9K0UR
98hzDKR9fvu6Vpk9UiphYvhb2cPlpg9i9amQDaPEPGe4Z3rcvJ1Eu8WyyHPu0xHj1BFwGq6H6S4s
bJY9pbdOokOc6ehCRpCS29EpOm/s/9HA1YUDVw88kEzcke/uU/+igrAHjQlWp/NRa/N8bH5sL5I/
XILmkhdykOdGXBoE3RV1e6pnkFoFYnmfVSw3yvF6FeJ6dNHaOQBLtuRKD5i03xhEJ2A1YuB6jqUW
odOjIZAz8yxBEsC/GIGqJT3iTqKQcy04ZH2G5JjdFIR3wQN69BGN1GedJTrIu2hAeRV0R0pRvLAk
7lnqhsL956K71oC9UPFYERXfxU3AlNoY4LDi966VaHNcvo5s1IYvNUkKvDq+Xje2yu9MZq9uIcxL
tc/yErDfEqHtdgtxRrDTbMIPs2nGKg6LSaLRlnngVHfsa/cVzesgAcMo/c2EUDoTagvAxWNOI76D
mPyf4sYupA7ZtUk9BwIOvoNrdFwfy3FbfJDzqb8yVVHDYqpDvv0ekLy/9ewGioTP9FG0kpATx5Zm
AMelv++uInY6pm+otrEV0QHBfHBSUD9+qNcnigeCDVmCU3eUGxfX+TazR9EqZDNUNV6TDlpsN3cV
1sj23pkVSrMeDz/5F90C+s/KptQ0rcpW7r+bPFvfno2sYs9OFJM15nUpsf0TTpDXk3cgF0y+xIlb
h8XtuaRLyvZAtGx9rFIRD4Wifk3f1YuOvam/yzXU8mB+KR25bMA4zA6Zn/GLNByWXuOVltGGh4O4
J/A+ZffQ5AupXb0DBSor3tY9IfM9afTGTS8ORiLFjtOdaqVC5DEMscndiUNLIx7YCVJQo4XXl8mN
0pwjcgbuGGVtPmcDab6VHJsSzOpY/5eip2h0ywY0mjg6JAKmB+9L1ti8+Iwy+YIq6dQ0HvjWq2i8
VBDUdZ9WSBaR5zpSnkmlr3IMOVmOTg7kpz4sIe/2cLT73Pc8ICuEiWQdnugaf8N2Iwqgm/uW1GlM
GSWWVTkYOyyAfjWYmtd139z+xy0VashC2RrNWVI73lSdz+ZJBXOSZoNh2ctwzxV2HbRvKlXAPVuz
qnuCNChgsRQePrDArkyApmppm0OuAO6lkIqHPDwZl/tNlmmjKfxMOKNmxg+JqFjBVnmhCWqj+aJq
UypjJ4g2qnksuwqB9jFvKPT/9DPsUviTxdtvNt3K/LPiJlsQyZ5tX6+yELjc/jkbQtLiyB2dgKRJ
ULgEIgMn76ZjiMumR4Dau+B/AmCD5G1w0nRfjGmwD+4GHjOUCNGfBwL5+2qsTC8h0u0nCUV6OFx1
7eEx1j5khEigzU704PwCGIiMhOb1BMe7U1D/iWfvHn2CinsMZA97ovhfTMjhYoou83hn5yMbeski
qoHCT+jUZsDFNuBcdrPg6rzplFFzAAYaT0D3kF77dutaJw1g6Ler3AYIwY7lNsbv4HoqiQpv6IM1
OzLkvC9twQC1J3Z+V8EwzJU6LOhsAkCPD5kFpe++/sfFoenebLwIuO/Nx2XktHS4xAKUczb7C0dP
1GmYn0GSZbqe4gihZ4Z5Tj6FdUJMK0IUXHWJKG2N7GbKJUpt+MAl8eq9eJ5ZwikIJm92aELDBTvO
O9xm1aj5bOmLg3/8qezu2yB9HTAHDULZPbcvVxUc9gHQf9mll7Xqtw58/87vhbd2PnNyP6vLDmew
vckdtf0ZuftyI3xulvZqhZGtZD2VLO5BvrmLQcxQGRiHCJWdq476ddCpQSJxyIoT/kwkAKfXrGPa
STAwRPXY9/wQzc5pMMVYxokWlbpq6GSNY/w3ODdyL9DpBO+PgzdbpNLys4ZEaUy7/CUIPn4pR2b5
7oWQTA+u9CGcx700IS05WkYRe54yFAT0oHTuKpaKr+yeW2+8MTqRxITgptDmvKzPuVFcdGRyCQnA
O6cqVPLzoznrtmxy5jDm5ZIXd93Q/yWD8hiRLNv5Pz+aJLmeKrzfs7igRM514o3A7UKi24WZWyOM
yQpufagrF2UJSs96txdflAoQWxXKjSfZ7TunAuEFD/4243kBGgLlPTCvykTYXAPbpNDCI8GC4Ez0
GpLYI67CEobhcZaRAdPr5o4cI+UTjLvhfEJoaGtoCVgm5LuK/9D0w+6sw8G7gn3fl+iUNB8/sLEe
N4seCGXcLI4xeTtSvMk5XOMnKu3U8aNAFTqf+N8dKsT4A/f+IO3hPFRVLii8ThLBTzB6CbBLruoT
Yp6rNLRmJRWo1lxR8B/F6LFaSSmOhee3QLxeJ11OdICOWChBAR+Q44aS5QWlyA/8+ME/VxNMVPjP
phuCfEw+y7H3Nn95RuySgO+gQXezG3ea6wUVA5FpK4ook5Z+iojcW/8ZNau+aBqxKzGVOEfUsWmV
1Ne27KW5M/MrOeKMeMDcQYYk2TnjeHK5c3mCl14Euwtb+QNO4cd5zlN+/U0BSWQg8QoZLLHtgbNK
c4zxHoVWchp4k1eeNqL7eBs65HWbl1kDCaF/8BWo/MQ6J3X0YFiz1z1OtSxbgkI0LzTPVe+3I/Zb
3Rnhf/xLub9qP5U/aw77xO6Gt79F+zyxXIzLtLrSULLm7uw4pRhZFFEhT/ScYlW/Pr8DxLqMEpPy
n8H/1GcH8EbP+CAyENs+gKxHLz80+7E84VWkiduE7fvhX4bZcPVbu4uh0gbGcG57t1tKWJDLToeh
ba3DFvF5SLGSqa0oy/znKRuRPjehtqzGYlU0DeW/fvXOICAVGVX8uXON1FdNEbrBshnNLg5/SAQe
0Tt6XUQ2v9JWQEypIXH1d8D5/y7lLQFYQQBrYv41JxDTxMR7/qD+T2bzz8kVdQ097iuzTY1xvg3y
gNGh7RUZxNsaoDarHzzCOPqVBEueoP+G04srcZ/d5dZDE0r72M6CYGwGn2msQL2eZhcB3RwcK+ai
ADVUxIQX43iXldpBurFaJgS0wLqDLFBB0gz04U/FcoXMRNxjgW7rDGy3c5GAUNhdhz1PWtA2v41y
WbH6K8ngZqVP3bVAL4s4Uegrg8PALVh8IpOQvjffgCHI67dX++85NgI76U6r0YNilCufy02XMq3k
PlcKngw7omZZuaoBIWsHXPLmJNqJTN+yJUiCztn1wA6U4QkwEttZXfiMZqUSMtEsAhg5hGa1BHAF
p1yYiM1iHzELe9y6PMFWeDdQ3p1rTx24CVu531Cli36T/xzW3zuA0nNbIEDgCMz0Wkb5XF+OKqiA
UYB2Fv43AIxC32B8Qs7QLmKDc38Sp8nt68QhwBVyGoL2FbebMl8u+64RYNSr/dBxh4tduNqCR3Ji
C9RWobVpJPKUsvNWRvV/dgiDRZ/wD7kgpUF9HMmQ88m0wbMgxYwoa+DWgW95z00/OcZlD3bGnmVX
IHdFhXdJ+GiJckmVVl4E3WUYOkc1vS1Wv/YgeTC7Z0sMpqHB4C+IhunI+DePIRoDQtRl+tHbmOA/
JzjOKVapNZrn0vcDopCGOa65F2UOH8Z+XPnS2EpqKFi3PhUyU0tJKJOkTCwoHFG6iQ7/f0ELtQ49
ylMOvZGHFqEYpci0Er64yQ6CT4eWxySryUCcoqaj0k4RT33E+pgRLPdSxhvtcv9vNQTRmr4Nci4i
HZ5pmUXW6uSvvBYguiOjiBWPV2LA3LAu99fZePzzIhWxEuWVuesuDPsTZYuEkzdW1ax9Ok1+6QmH
j56V9ENIGJDQSZvVtHKQKpcPcBdNbaxBlwNSTYOypVoyPsDbf2x2jCtWIEccyZ0Bk3lfVr/EoevD
/8wlMfAOSB1mMTBMMvDh4X9DM1SaNSpWjWHjpgUQGOwMrHWjxjsdPlNqaqH7O/hseLK4WArlLD15
EBPwX3DUujaqge3K8aVhnt4ettQmjg6SFSvvCSHdIFRl4qeIPD3mmo7ipTyIa7ph2xfDVUZrEVyj
T+Vrh5mLQzsQNJCy7bl5JCHN907ejSSw6S2g92gEyhaTFeEne9tEnCkfe2ZPmZxGI47ywO5PpJ0X
AVc5yJtmrCa8MJbgRtbxp6rR2Swx12VbWloRMOzAfynz6y7/NNq9R76kqkGUygpkoEtdQ44NfVJR
EkCORhq198nWekPgrEj3XBcoHq7Vl0guAJhXTaxTWr8xbWdVWVbkTk5VWeK/KGRiPx55zBXZazSI
vkOoz7KuevhFViVaEjAeD9k5rLG/cJctrjacxLu6cUzgaFPGESXXZC0I0aqZa0ndAWhNp/Xa59o8
d3qCwPobT/za+bHmmKgE7S+ugyquLHH2N9KTUPcb8F2NATtOftFXzjUU/i8XEXiQoeyX2IOXr2KH
qnv3PQMg+MLAp9JH5dizMJqZcqYlE6gjgrtj9nC7tVvVtR8DN/KfdZer6TqG0d46WHtrj5NVax+9
xMgb+d/r8nJLv7bU39DfsKaXKf+C4FunUx8ExoBITsua53OtiBo4u5PkNKuMSfO3ys9eCCnj9T3a
xO912sCL6UksAku+43A63SZlYNo3yfxs6HWR2zs3esf8QaSHeeySS4ITp0rq8n49KyVovNzplrHf
BIB9QwZ27sKZuZXozql8TA8cyqSfd4P4dIdnDLeKxpntAdf/rIB8QzceRZ0P7MJD3wHwgkgwoYTU
bmU3L/OkSckred+Sc8JZSR4LIUzc4N0/5tVblKYE6uoFqErmKoAgXu27MMcNn+4xrTU65p69xzFw
jwDtG1kUNxGO/J06bvID6oQ3DfaoV6aN4VP8+InZFco1O0aicVDLyZIN+N7FPu4XtSiqP6Y42P62
xWFZAHq10W4AhYgpx6UrRHwzqn0PoNPlrumDZa0F0kazfl+PUyW1MFM33mA75tMPjVDTBU33DDgR
U6041HH5UCMPAFGFmpWOWslBq+k2yQ8RgZ3bViURBP15mhrS0jgik9AMlkln8BtSz6NqLBfTSFO3
cUZJL/zK5XtC9RA+L6bz9ifdo+88b6drKrOYkBw/VGGdEm87DWHjbBu+ncZ2fuwcTN/rOmf8IRJz
aUfUYmug1+Crgj7TO9GNKdxa7pCljo38gKqaA/hSWkFSIN6qs7WzqO9tBww7F05xCCLIXRw6Dcty
JGSV/W3asNn4dE9uTFyrKURcTv1RhIta0LeBKmio4K06UbmeLRzbUConoVXOoGRrlK33PLvDgk9U
4KB7/VgRdLb8mjt0YocnkK9y/q6sNQwJEdsr+NjRYe305vcGIxzruypI3P/O7UzyP9I0QxJsXith
+3OlQ8oYXgvDdVjvn7qIZSpRITiOorBNgSK7NEC4Uk9oS1GvNxF6QAZixGFwahy9h6EHLb3yQ4xM
xQwNEqLmWmOXI2Zj1saY2PT7H5EqhQrMv2wGmILIOiaLA/Iwtwane+nd4dvGa4r2IMUjSHbEA9wu
rKdBvfX72GqDoLpNRI3R9GL3UNOvEqrFOqekD4Yb/WE1bJAUfnfVyeItDBsv5xQ+dW8q7u9mMIkX
ZTY5HMnhgT8gJkHczuG6NF18zPk2+j/X1+VPMttiDkBOR9E+cXPgRkpg0mXQegCn1n6kxs78dIFo
uOR5J9PBIwQs/0v2xbPQteN92oY73B22N5yp0Dm4iMgf41XCMdU+0vPWYNEEPdJMfoIRQYhxEAbC
ovIbDf990doOJY0y5oCdzSRyupg0K15eaTSVdqb4MjpwuB/uIUmoMIyaugSp3/LVZCsfZwytQGmb
vHkroluT6eadI9um2cpWahIgNLpVEwOUFAHAOlk/OmHj5npDqjjlHfrDjjYV67KVCJ6dHOygtiC7
ayIz1zLUMwUGV+f2JEdbp73oI8PdKP5UfqwtRf7yVwHsg3cf8AzD519vJjI/sHBVOgKEhqA5+DQQ
cjyO2YvagVVTp9+PfU475ynbVSie/ckkySYZDPuzKekaXTvdjFFOYWpMTsixJdlRyUD2n80Kh7gy
fzcnag+OVzTW+AR6b8zmVISNeiiqaQre+KY7HG/JfWPkYTRfu7xBEf36Oas4is/ZwX/JM1r8dQ1R
lJ4K71WK7hAADGa/hZeN9hZqvYJOlFgM9zoaIESnUy9tIR6ccK4EQqGVcDRBoJxabD0EEhJ7VLfC
XLIX9illZ9gkVD2yIBASH2Wssg37FKk2L2Xm+anwb6OzOXHVqtQoSoa0MT4URj0uWTSe9nE8godv
6d5SBFlY5iVf5/aF9VcQ37pa2F3z/nNtyRVOUe9G9FkfJRrw3T89k3cvL5hkQwoK00E599WO1XF5
9Eg3fip3q9TRuyhcxs/WE9oZvvV16y6W1hzkjpV5eDYBfa8eGfoV7V8dSgw4VIc/5dve//f+UTP8
Qz8j59u/wR66W27DKcgqtPbDWSoWxfq8Uk68TdPUKbvog8Jna+aJQFaVYyRvfWnDQVYKOr8f6/Mv
Zp/i4s5k3yqEBgkhhya6QgQaoHaot5GZ6qzVXxr442tXMmJx37/N40i+prTdEULwL3Gb4RH07VVV
h3vNMj68P1V1lj+LyaJtyPrf9K8ZbBi1Zd+T3iRokJ40ApnIpZKK0m8vacPB3L/URFvERynf4BrG
hIo+yXMYd/odGx4WrFmWI2MUhuN7nckRXwIVCe+NW4h2xqw3D7tm3JIO/cIFyib7mfMW6ztyS9BA
I8q0lRQFrk/TZxtxificYaY3g56SGKD3VrcNqSHldN4crv3Hya1aOzwt8juIs5LckGs09qRgxYJp
AnLmAYVPB8OBwiRzsw7mtfmobZ3shkl4WcDjkfQ90JasMSt3H2BrxBVMFfL6pEqZgK6slBaxs4hw
y/ZmAm8AnoXHYtLTYbYBqDi63g4ciXBw3CsYsaFGN9VyApgUV5hH2tz4nGI2RKorG1ha8uyUxrfd
+YyKJ9nN3HISHIqkMJ1njpR+xCJ7P1YDp8EOWS9Dubv5twqfYOZyD3FJCo+1jDX7hZP7GM+6DjeJ
UzsFUBTVYYP8w6X9T4QDgQ+GohTc7yPfc8KxsTVIftSOB/cMnFt4uG6D9CFB0OWSinGvMpgsLNB9
g1gXaCJZczp+r6LTNrD0Vz+BjuAbJwRigIuilPujn/sEI28SrMA8yXahNC1oFtCwfZviXNX92u3P
8rilMh1VEV8WFkhICO0XBhG0HpVV5iVp0CylF4CkDQPxBs1ka3RWRJ6EUQ0B4CD4SOVKQSjBQnZc
O4TRwcvABhYSln1b94S5K6oGKkah6KF/HerVV4uGk9o85BGhkVVZBVYdLGxaiC1x+fsSWoFDXCeR
sdx2dEooTYx4I4zFdLfKCwf8Dwrm2wY/Fcgva87jRGKvvHTp6Ta2NTzYmKM4G4RUycg2sJ6YvbRs
7bGelmboRmlSTCsXQOP3POal5O1DUbI8EPzzvEIJIStqgcg07kiyLS5SGRJOfEQpSmMhUW7tH8Ef
4DfvZTA6MxrYZ/6C75iLNCI8Y79ETs4XD0L8WsAiUDas6Q5pcBjIn/PMBjLoPhyR9rTKy2BZaoUy
WpYnjtJ0As6j6+17G5RGWdE/WsBsWdObc/plM+5uAaRo0i1UvW+8c7W2CNmdEeMvmyZOlgj4QOLF
tx1c1n8AaKUDTZ0mjSrPDktFqXhixcSy71LQxjSoIryMfazRWWK45D3Uxhrfl0j4K/knS4VEa25H
FPMBxCrz4c3ODpL6DdHDpDvFMyWLU0TWb0LaITFDCAsqIgaYRAzSutjFBHQh4nGdxbyytEs6XL+i
KtVpbHyfRicaigW/IGfMb6ukdvUzQ20XU7AJ2MLyddACUNZxBrjqOovyXLwXsApgCyB0Dj5N/1WY
Yzsl413KhPYws6mQxf+IEMINJ4EWo62uxNQgY0WLFYh5F2nh2V0D9VsPdmG02qbpvs3GNYTuQSl0
bTbZXaV1WKbOmh058vm3z04/AomzniruJa3iEPolMOBTTCvsHa7Y2h9FrNwt+AQdqC5qrX2Bh6Dn
bmmNn/Ec5DywPPWngZ62bOILVzslfa3QMpICMjv5NyXuY2z64x/GTOLQ82cXcqPsweAb+SOjKbUt
8SdLZz7Knv7BFZt6za6CpxZ73q0n0ZEA56Qa8uNlsc6c+j20xMILtsbKqUpBNMPx96JjE9gFFeGr
CGNcTbb6R70FF5gF5B+1hYRn3zvZP7w9w5iymWkkXarnrden6kDlx/xKeMT+GK1ou51H9Gx4YLVP
q2XF5goC4stE7NmPrV18rhylyq35cdHS9zTN5aGHoHDaKHcK/9dBd8uw7YS2OoeO9VqTqXbMwiz3
RUK3nUdWzEshYPlwbj+G95apI3eJjT4xMceOCLwekMcQnC+/RSvdOlUE8nXiGbfi2WBcXffZwp6+
PeYqukWSqVEkizlGdU5rCEilVCvTkxV9CVFVSkAE9lzZXCEzpfr0Nmog+WCJVpEOsX4OfYvUkm7m
5yZ0m28yMEOrTlNE0hjYRwETptscU+ZK7DAY3oWVEz2wgW7WX7ZlVe+biqYfpz5EF4YCzEDa7xAF
CYpgMSSphZCehQsIOMumHwhhrRT0tqm4mj9vg+Trk9+y5aNNKyywvJzzeKOz2cgA09GFIwiDqrFS
vwj7+29xJNazCisc+/bc14Dsl3qYSYAnkbi+YstUXzuBhfwBfdlFKA31FwBovtuEn50WGO+IwaGz
tIQOy5029cwROj7jgap5H07oEfFdqfKhWfHHEwhD78PCXaNavbfOEcJjKRgT80VEtuHze3Eg5i5b
V4di3s7AoNBzQRrWlIVumfMJkesrLusPObhNMTUK2yM+YnIqoKO5DwRgrI+J4O+DRB0aBZIqNZbb
SECK+29UxEX8lwK/JDwkvninHNkBGqxo6m2mjemAj16zoAkEXwXtSjFuqvy2Yj/0J+hc85dxfsnm
JhDp8o7DaFhjtuj4KAkhBDq1yLMz641XJkxbYJ0VT8y3G9QLyYEcfTLT98A2jU8Bgdg/j5bn6fZe
Rt+5y90fZurQn3iJ9uUCG736916h3tVtoUGqMJnAXbk9h3OeiBuNstKEJx4kXZgjh+WpIrCBcfhE
DuUV8XTnYHVPH3TDcPyJw/KMSj5bIXPpJ2Qey5/ui2OugioEVb1dB1l5sm3dspUYma8Bps8ZLMQZ
hxCjz5fUQu/cPTWDof42m/SvnuZ+ixsdz9U4duf7ldL+6stGKc1ePrdovFZ0pHLIndQgicQkci0c
0XspaDNOjMOavS52bsu4aV4t9pmmBNIKfEYv8kkt32z6zwmUlejhFAihbAohECMYVtRP3vuo5+Lj
EPSPFI/IMJb+OYAUyHDs5ELdhDIFenQHiZpUGyHlWW8tcW6GRYf7O3aoqnV3QMtUfhf/UkAdNzrH
YdDHkFOMHmdiQWKpFZ5wmkI9jj6hz6pVQ17HLJxPTreF0juszIoQo8hjh6wvhwGMhTNv3UNRSL4b
zAYxNwDhMox1FyqLHgg67vFNxge18llVBv0s3fT0KsR0h4NApN7AyxQQUugA27jvWxLjwOeWJHQN
tL4LnJ3Q5BvfNhVsi3jFeTj1zVWm7Pc0hS0qJUdn7aWzqfEcY5B3KxtLfyBjK9wi5yr2xM7dNmf0
1GK2I5rQaYRa6gec0B+wjC7DCTeSlJgJz50V+w6ZwsgW2xlS2H1I6A/pdw5YPFIhtkUlg/9NEntp
LL5GxLtTw8GprISYyjFqp7c4JRgF3LmniBa1KVTARwRHe8JqJOmsPtLOJ9X9TOldaF6x7cb/2gkR
E6UDYkrpstxXUdZfoAPuVEhWvsrIOYKy1NbDXiUv1ZsmJd10/mAEiYX3bdJZSiyTmbDBhI4JQlrF
VreatbMgEdGhz9cwtHJ9ptviKSJ0fKF4svv2Tw//vrQHR+cANqHxrrQNPOgLZA+swyLSWKKemaE6
stWdtiw9vde6g9OYNnopwp+iAHPvX6c6ZnOm4t75ENavigrJGs415stKFtrYUzIXtbCsveOcBEaM
TcyC6g1+ZKdDH/xa2lQyIdxmt3fUR7rDj6P5VayuN9jOIHQ6kiGX7QSLuGZ4L7az7OpPgUu+o8jW
So31j0SGOg67P8bKAb/Z0dpb+6T2sTapjZ9XIRUmc3D66MuTqgaE95uJBce9yw1m4ipyX+0Vi0ep
yCt1BthvNdLoxyEIvuu+IJIjC30Q/Z8l+E+UYw567hfcE9QckzrUn766SlgNC9swwpvwVeVRq8dp
V+jyh3wT2XTAxTltsCDLhYnC1d4cGuob1AngWPrMh2Zf02Byufu/WR0E4pboUPA+tRfozAbHaw5/
wXL0dcYJxrcV9cR+4oG5ZmPrA/7jOdqL9Qg6wky4le4vLCCrhxk/ZUmmHcLR5HgfvaP2tiDDq66b
ZtnKn3s4GRKwRYIg75XQmQ0dPbpTblrO5/eGu3lSFWebKpe8O65DN6J1mYVl36BF0oD3x0qU1BuT
vBZrLTN8l7UrQ9AmpdrP2+FZ23OGT3vAxJOnU3hLM2CQKX4lPHkzmjOJIoT/v9AmHUXFZkh4vNur
URO24fTWHAGjJzWJIqXDIKiRP5rRMCf585bQG8UU8Wuod3sZ5tKLwDqj/CcvuzNxZWw1VDLSwSaz
uixUm/SRNUuf8wxH2igcui7JFCK+owCneHCvINkNjs5HSWjRi9qewDsc6SGDsY9x0+nsxd4WhbwV
JLxDte3poHaiogUhmYe+x5fC2yOHglG9MNCR3mzFCuxyWlK3MIgQuEdkMSteIAd/qSIVtbS6v47a
CIAMWV7xtmctvoJOSdByZruUzIa1LnN9qoMgSDBAJkWzk6Y3NFumJfVup7SJ8lzzD6WFpT+2mPSW
3cpbzBD0R5Z2H3lsSLHcQoUSXss6MoHqDGo9vbA3zQR2IT+lN5FR7heZgxkv0XarfJouFWFRNvdl
K0dLeF2ph/SejaOrLsq5DF66NmeabnuxnYv1sonaWv5MMH1RQAigBbb3gWNPf1PCQRaq1TyV3n0F
R22i+ka/dzAqIOsbGYJcqlBEJWFNp7m/a6Od+mLdysQW1RLsJh8/lwypmBdhQhm1nIqh0t1u0OX4
UsyVw0VyGfszELWi3Bmj206lRmecwyhSi8Tsi99aMxB329Qkfw/hPt9NEBJ0nFOWO4aQLK4Vxyyd
g42C+gJ062bMdcXqRAkydBb6tn9Lnb9OyG6paru9R68HjSvuVLA3vTaGVb4IpDrPQVPU4hmy7c91
kDiDBpkTnCD2sba8bpfsKyB0hQavDmToXjpi6HP9thUfNgJ+O1Ia/gyatKeL9tbAJGqxLXv02W5f
hV3T6FtNf3Ps+QUsC+fSAsV0EQK+XcwhUIWLl1FJEQYUJuXdke4rgqHbyTzbHywoj4UoBydANjOX
n3EAWjILlnYAa2EcS8Q+vdk+uDqMFZqTfVQOX7FBsw/dzjnF0ovzg/WKPHagay4wIhdlz+qV4o+k
euXmRqOozrjMFykGxj6R6qze03fA2Fu22EogHzHZB6Zh0Kg8yWFbPbllkBSLvjPZeA62ynf6Flmt
ehqLLeM98/1VsGYSmC3VgffxKHQGAa5CtkqjSwfGC3MiuwPz3+UVoAjv0s8iVGhX/yGM5cdL4kgl
Gv/r40VUujhbUs93e1wNPC1SiEbdPslibllpu01+p8ZDLEb2pqrlw7XY7yICYr8qnsr29k0aoPSC
N8gWg8CM7o9LeJSl8xcGQ7hzZE2aOKwtrrDJ0DRi4xW3119G69IcPYoRrf1qdgNlMZ8SMKGL6sHX
yZ1UwTIAgpttbRSLLlFhejoAGwWLlxMr0IwQ1CFkVKNyujFPYfyMtH10te+86Fo7yc1wgxptMDqf
QuPdwyM6cgFRko8d4uTIM1LNZ52yJ0zQywmpcbPPD42qpLwvakoytQbKPvP0/Nr6mDoKfn44VVDr
mC43aHVICxyPtK2cwPgTNgyKe+ndwuuSYh4SQbPxpc3VhUu3fLQwl5+iMDqyhelmbU2iwYRgsAPT
7413L7IVeLrjd49WmqWvJ3C9QnIgkcEJOhaZU9aaMfS5STnjJ8gHuD7mfGt34mUGdR1utM5VrXjS
mZQmlq2QnEtJzbdOjRPqowmz4Q9hmA4e7kO2yjY4FhSzLkjefwmUuUh36IGi/4pkcZVZfPGLih+p
zB8xuWBRxtiOExj6oy36HYUMl2RtTtwiGxIF0inVEPqOdAAY+OB0JhGyBT+pBINVrYJp8g9zcEoF
PqQLhq5Hxkni6ZLQWQgR4IbUSJH/mBT5FAR7WekPSkMoomgTUrkLHvS8ymy867sNoeK6cod4hKnO
/mvnKCl7a4r8C4hZlKFirCbGmxQhJwUGlU3HBaiariteVUFTDjjJyYL6RMsQbF8GuDNG2oh8ZOy3
ZVITKj2j3AoDCCxw0cVuQVcijd8Leep6QUgA9Ie+Ia/qU7l3+rV3exhZMtuo43vmQN+3MWX3qSWR
Hn2+9CVXWyytAfkZjZDCuj+K8cPyjnYvvFIwVmn/ZQjL8hkhHBaArCXxMgg7L7I15KlIAUclsCrR
7/+Ol4O1Uw2Gl0VYxsrw3Ibrgn9JRCHvJNpP2CMIyPyhV4yaD/RUbaIIjFvD4Zd8o9ZMhLrg4Slu
FQFAIUJ0ZcTInveqm0Ecg2Q30o6dWmNhFalPiP9lrx0cmnVoTuBjPE6ySlq+v6sV8tXPZapzIBcX
a10bEcrWnLjgP78DdmggJWzOYkrKndelwj0sg2UAf9n81Th36N+Dvv0CFxrG2QiUm5IuJxVYoT4J
J+Rzy8R9G2Q3JWnWGhV2dq9wr1qgKWC7L9xFdUyDJ4BUgGOwKzC3CiTMqK7K/3tdQRppwEP3IiNB
S++nPwemmMyKEAfdaGqg6aipNOXYhB2olhLPqIYP2kG5UPpjKffGwv4hccqreG3PMbrZeqr8/HW1
OmmghUVTXeN8ufslJRXCAy0csDqFYWcdnmu6g8v784qirvL7sp4YSQR6IHgjbdOBkOlHVGGJRCOk
wPWbbI/XTRm2hXmFFxnIQbhZujmBwjFvToX5TMwgbVFiA9a6fPZySbi5TVsAVeJHQaQD63RHiOp/
PwRmHzpq48gWRh8fL6T74wSWTTDDheYYCL/vyYJxZPaZG5+Cg/4i/vFxh+r7xgvT65mTpKyX4Cbx
7Kl9EKyS0Hl94OWpmrd3IY47vAgnG8KBdPRvdIf1pfnuc3J3QKc9vSms+w9wwX6cpGpBnYi6CB3m
zsj5i2qOzddOjmj9I4fmWija4fYkZ4oOE6vEsOXKu7wXU4IsmctTAyJLj74afpndGADphv+duMTo
gBLe5MriKrCi7jNjcwl7lxU1tyg0LLvN3MbXXzyj9aiKs6Q5q0rYJyu/Kp/vJ5oPdE/Ru36G2kLt
QK5IODPPNGG65ax+UFBOps/gb1NzQqjs0zg3RkM29cK8ZSKOGjEUz/Kqvo5IYXl1KFzwubBseDF6
QQ1fZR5/VmFFgXOdMd08Bf3u6NtDr+OnUyjS+EmK/v3/kWrtPD6CoLADoI1rZmMC20BJpmcHrcpx
cjuTq+nU0AMztCfhyfBvXqIOFXc5tQ/IarWvtxhwOwjwVWJQeNNPPTPkwn5Am8eooEu4GPYsYzCY
j9eD6dU5ZdJkYQ61G0Snk8EXSMAMRsY+7T6IjmJX01TrhRqpCUdyom+PdhVfMsazRZTyukq1WRfF
hDTFf9pBYmD0NDSpJEJ6BsPN4uz0oXMavvkqleLwqlDbr1UshYkUs4HWaHoyN616OK8f2usAtJs5
2+v8RRNep8K5bY9LBBe/upCa6ZRkXx1+7VdEc16ruaNT0s3yjc1dIxk3RzYySnSx/Utpt1+5q6Zf
QIPxeLZoLnFbeRhXefgEzL6xdAFlgU92he97RT5K21F1gRFn8ytfnIUuF1xyYtHEUsfT8C9pAxCT
sHZoYlNcZWVVlJHkW7jnERCR9fay4Jjkqp957qdFOaT5XmIJ/mHLzayK+KqikmcltjLiQ/4pORbL
OR0IayReZczuLcDnsT/rWVUpq4Yjw/TJYUJIp69dAjWW31Eivux05yakBMVpqURyE5Ahou6AViZm
HL7+4iQ1np8ficl6NUgnxjpKSInAsXksvRgUWizIb20D/8nwWyvNBfL11UUerTuh7ePGkJKN50Z+
m7u+UhMbjtdbCW4RjGoMsypA1E63a3+/7uYAgNsdzLo+UqGZYs2lTt9+DYJJWIyNedsLWeX6ffMc
RIwwt0cf98vkBpEacOafrBU+I6dieBSOQseCww1AXpMFz4uXWwVEgyKGWqCb8rlYVnu7tp8wxu/9
nrJu1IQOaAvA1c6QVVFtBZ3Y2HDoEJXz8GIQzq/nhalC2rPFpnY18GxwPl9SS312qz5101qNvrCd
c22ku7/hQjzRZf/QmdDrNskh6TtJemkqdMNNN7aMSxoWNLUOcciEE6YYPJEcH4qxfdwniy4EMfmt
wLxJ5YAMmmx2llbIcE8OOqQkC2AYqP/tVOkwAXHEqgJ0cLTeVS9D5I7BYg4fWdIK504axce4zuah
87RphvBOlI1LVcho8PNK1PjPPeiOfCXZDTKXvanigp7jxSv69r1laJJHTU1FqBJPJcmKa0HzqLyK
r6/LWWYuh0bP+gXRr+ywhI44gW7Yf+epp1R22f7Tm5Tnoph5ZpRzFt10hk3hT1LXU05ebUYZ41+X
GYCda+D2VmBxFR9FVgJSwYeDf2Xu8WnaEaaAsatQWQNzwIY6AbOwerh+Gsqpt0oUU+qaUesLScMj
jBPBCYIewMCTE5X2/r1ar5kS+y5r0tAt+bQNDdbJNbCJexLBLRn8iHiGT9F5wpzUdEzqznGqXp2a
L8mSG7ZKyXiEaoFINZ2ug6g9C5o7T5KnDKz5KY1s9EwjKCBSCZyU/ZnKZG49uyCwkows7OFdHO4O
kRj7IW3lIA89kWRw/6kLgQUoc2cCsq+ZEGx+MGYWKazchm3DDatX2gC39RArmstmJ0CjEpl4aq/+
exvXA0NTpftlaa64DexTh7Rid7byKK6wEtfmiHxR26mbnMnZc4+XOi3VCHKlT83zoHMvo6gZtZS3
GKoe6B7i1VcsMYMvf4OfDogxDps23+vEq1vzPRs18D+zlAx4Atx7tHXnN2vfalhgGmK0/AfDMK8n
VWw9r5wAtXs5/cEKR52YWsdnccagfyNUpP7gNEC6Du2QUfvDYU9fSYp0tmVh0rcLzLdHq+EshwuD
yr6uV7c50vdPbGhvlqdQn4mlx1f0TWIT5IkUZOg9k5dK4xjgmKybsqGB7Q3M+A2FaUEGXL+v1PLK
lXvL8DzDYbkhxwGatsE0ATWqV0qyYiDuY2aM5U/Rpsa+qXeBnYDdyE3Jk9Cz0s4nRw9n8lex2aMb
BsCEwm7GltI3pdeLexo7tcVrbgYGfhmMm8CHacQkkxZAAmCvwgQp965Mqs0ka+bg5zAYaW46x0U2
J2FGiM+URnCny9C7MFQyUxWB7kj5ptqKEhY6RaKqdxuhn6mlYe4IFYaB5nzSt1wa3z4uHdC0HZlL
UXXkVBjRB0wBa+KMyB5MbF6DdrWD3TXspL4UZdAmZ7rxqfyxOn+0XCpGSvLalrT07aM/O3qv+ZbJ
4PPA2pAJ4jNmvRaLmIMi2gQvOXt3xXuvPD2h5z+B24dJqPJE6CA78Hk+RxK//Ai+yunzVN3V8N5V
hgzrCpf/yuuGj2MtnaacQMQmhZ8XM8bqzd2LzqRt848W3lUnafPpoCFyx0D65rQBZWiGq8xSGDNh
Fc70R9jfPoM7zJ8kr39jmZ1VDRfrc64nXBkhHzTNyV6DEGpPfevY3PBdVqUHi2X0VLxAfrOrabPY
mhvJi2v0NU7Jsf2ab9Riu8Gm1vU8pJi/afCwtSLZm7ag2xc8SQe9t2it1BywPSk/capgJLgcK7i1
Siowk137eGsIqAzzvF92cANQib/qpncWLNoitbj5hEWuVj+9zy/Q2VMK9hj3hUwccqVFEJV32DvH
N+hXGVI+Qg1v4FrH4WskRoEZgY2mryQiCA5aAP1ZHWIpkydaeFGS6ttG9pMY9twuYwYl3cH+affQ
PRvMWuuRvtFblBtTDt/iQrDmogOGQIRYLNHluVIY+DBoCdp//AyjbL+O9qYK0HjtpbIPBlB30SWn
/10CFUn3Y2LqdVmvBj5z0JH+4msflmYNBIQhPG1uUs2D8EMKLvL8e5C5QKMxWlyzA4wZagVzzW5c
OX7DA+otZEKqlz8ORe6CoiDVZnZPlBvLUh05PeXz/hnUTz1cP0UBn4YwXrNtbe8dFr1sQYTnRGDh
vjv8W7Uj5P/4OWSatwQclUue8MKS4G1ELEjCMbLWoJGF3sjoEQDRtsswPfD/pnn5GML8dVvtCq4M
2m1iLUM3/0x5zVEdc3Hp61SSWQHcaE6edksnEa8Bdjkjxwi3zxgTxVBw+WmidozFvdNzvp0PixBj
lazODQG2IlRc1WzsEDl1XjYKbN+J1l2v20sjgg+z5MVn45QPTNoqIcOkuV7ayyPnjPmL70NrMrXt
DV6zmaKtSPKGCoF+Y/k3GCcZ+rK8y1pTXd897diR5R7/+KkDKFnjHGjsOcHP+oK7mgYxBsylpfie
9PFKIWK9A6C2ghszvFELLXjnQSY+LFcRUQjfDzltizabYC3kSVoY/6BWJXGdnLHDyOMz4Zxmsjz9
swGQKB+SB7zzk096RPlgeKtsBRzOXaRctPurtPGqLE/RqJfczMZuPKJ0iHuhAICT1tLT6qF3shnM
6o6eRaDld7RYP4IrjG/AQZALNB0EO2Q95hRzZ5/Lfr7/yW6pIfrMeQWaSpEl4ODkVFg1poWo4zy8
PLhjzmePXYNdL58wXm0JyVlcKC7ocpKKkoysSXT7JZS4rw50mv65wXA/cMm8FsSiJdOKrTmPbIQh
CUn+dAo/wdcopqGu6xee5O4U7+xgmYPbG5SdW+Tb0YHav6YDTTTQjmWFLskjH6ZomyNQkBEBhzWQ
xHO5tayp9YCc4ctU4q6SDcD4D1A6gmeKIBPc81zddF+4G/iIYvBuW/fXmfO018LZqwZU5BDSElDv
kB+iC1SlPfirqTle5valquPuVtcX4vCCF5+9M/mLDJrbhInlLOERL672iMpZIZO3VL3Eg0Lzfem+
tIGwN0l8sTe+ELNc+cBqODrZn5v+WTVls1f3XbySl9/57VtnRelyGXHfGkoOsNjOuoxCNeUP9ncZ
/RJNU9c7ULmvQzPN8tq56oxVtYJaUwOFe2p2YibI02SW0eY84Ozrx5Sq3qLCl6AEBlcX6qmBCOb8
wjmuSSF4V8/INJ5I6XwhPpad54q2+cr9mjZCso1G25J+/CLXoFCFCH3K/z104BcBVJxxgYopkpLf
F3lyg2+5aODbwAuJdYV86i9yDZbvkRRNYTldD6IkOgvt7CdiT++6/b6eFOjwZk4QtW+8H1rY4c5X
vTteAteX2j+FFJH82qha6hXm7PajPXrGqE180lMg64QKaJ5+y2VUTD8uDA/gsGaHKcvJqUF42BMl
XuObMbUEM2ojewdf4c+OnnjlhIEy51se+d5UQ9GPyQ/f1mVZMDOqwjn0QawP1INqYJ1gghq2lznQ
0GaSG1vqbVDt16G40/HY9nDYR1031K/OrOJ3mAXD4dU4TxKP7l1m2VjUJPJdYRe6cnwbjrcZV6b5
36/HZKrDp7lH8JPpTbBpHdpKDNi5TPsGzoEyeFugXI9QdizRLpULnuFX1FFTic/bFo9M1b8X/GNn
E4e4lKCGQQbrXdr9o+TPrLkRz3nYVcwOxW2QD5sJxo4p40CCGJ+/nTtJS9Y26wisG9syIzLjkMVZ
bOTDVFopCTO3+A/sopb7FZKxhaySItSVXXwK2RsT3Wil/mvYSBwYGXwsoe6tThcgYD1AL+FKXmgO
GYZ3N3/+Jmg/jyjiZXBzVOJ5snJKcw12GazXZ7tZpd/lGF2IBZetOCGMl/hQv5r4g2KpDUZT/8GD
+EcJ7Hwlbt2ZZ7qSpTJfFzjZ9bgFMwyafBilGq5hu3jHSWzT26kxTW4CZjSBwcs3PZEq5SCoOlvy
9m3Qsfb57MXU1BvTn+gx1HW82aFsMohYLzrNmvNBCFfPNnODBadJ3JnbVxbh+RixRbjKbUS4RGB2
aC2HLl2L9+2l4AXkpDJPZc+4wNmGCEMtEEcOSAxjxOUbFMcvbGaTHzFE+Lo1dbsKIy2aZ293XHla
YPljwB0tddE2xFJgKL0nVfjtoT4grp9/6vN1/pjVqNbKa9jsJ7uNKs/K2LvOx5DHCT0yoQpuGfgY
+xQCYVslNwdLp3AiqzCRoI4IihZMPQwCK1Ep6zoGz19iY1RjH9L3V6qQ43a7XZg+U+xZ9cYhau7y
TyNPXpAALiW6Ce3hhWIxaWMgCUnLSL2NhBA9M/fLr9L4nN4HHrawKb4mbzXJoePhPwGzOjVWS47w
wNJqISgdzUmxPnJp5f2BrYJYBVeJ9sBxGs2Pe6ue4vRMeAyWI/V2n61KTvPUtuNmpl+itM1ZWF06
DjDfgAkjDHJ05OTqX0itHbKW30v0AUk99lqy9bXlXEHnLjpk4Y34u0NGG6WPS5ivPVFvOMjsKeqt
cBmOBRCzVy9R6qDXCQ2fusZmLXC9OWwbmMOCsHlGYax2hQh5UWbnbhPFNTBBkxk/Whf9uJRhovEr
ooiHYLYDZxwP/zENd9+y+nNtz2aoLyc2DIFi46MCjz08y2FtJka0WPi/kDmD4Y92rT4nP/nbhwaJ
r2C2AWOYmWCKWQatpcLhWC05G6g1njF4WNoPYKnVmv5kErB/tQLAwKXVBbl1coUmpuWViBQXkmz0
s3KDOhrC9LOrmMR4A2vmrnZbQGGaxUcTG3gdHytrOq+qtMWazMTmRlbhLEmXmb36w7Vlt2AdTtOq
l/S9IO+MZgwAUkJb2fWTh/TK9DlmpFz5c7b5Hbv8l1RHYd8hrp8aQXGmCX6bKXei/OC3Xb8gFLMU
ZotQFYdgAucXnM+xYfEuS8KPgtm3M7uGR4VRc5yzZIfiIOsCe5r0Zb0UmaVq5+hcfzeQQJ9t4Sy3
kF2rV1fZq7rneI/VywXgqF4qQhEZvcdq1MpiWTe850LfCqXMMfNTSMy3KHq5SKdmhh/4eZKvTYNg
XXV8WY3Ov+O0aAbfTuwQ9U+04wYr0ksdXp54/OtpMm3z5f6Dwd5mgGUKVgAT6YozB4pSi47SyfOp
MPUu7Ia3hMzUNpXHy29xVrKE5Gj9nCAMDrTeG0r+rj5BV6JyzB/XGu+5M5e4ymRYKNve1vWcyDSg
40sMCQmS/TOER52pivcN4YTOfrVGqYp8lAjKCo04ho/zc1Ee/9qqJNqeW9RAcJLdtFI/BU9cJYi2
ZkqX1sbhnWU7PrszRa8OsBgEKsSgMEDrh4i3sZuaxYOPW/wjM3SFeXsC5aZ1lGedyObrjGVBv5aC
GdLOOWjzqqPDDNEecSHYec3NQnxPAR/JzkBGKpHsRX7Rb7CMAiSlIU0JsV2Ut29mmsrKPZdy0edW
rzBmj3zFSJSb6u49Ag1E7Qj+GBZjNJNDgPCZjLgFPjuAJh2OWUfHIbTW1ysOg8mUNND1nVVwMaHL
TmJGwWucV/mSXRkp/AbZC6XM0asEmXcveW0L2nUNE+xkYw3SlCiXcz4yaTFEgPHNOvIWjbmdRvWN
OdNGeIzRWynFuyZCej7WdD/Z+7qEyM/TZeVznEtzP88Rr9DfX285D71DgWOf1uYeY8fAuiONPo2D
ZXxI5B3RKkZUQSkO1HpovoPM6dheWmzzE98ZNqyfQIZoJ12XC8niAuPhywtj3dV2mx6/DJQ/cKNn
D1eoZ5lEPNtzzp6Ax0bUosoq3DLR8Q5kgCL4xPwzdWSKWiNfbSzUrsESrLE99e5ljJccEDbXd5OG
0Mo/4XcyNNMyctvs/lH8YhfuOII1uamZaFEJOB3yLRVdFbJKFfmGGNiEZp1crqznSsrU+vyfgvXq
s8CUFikslEL5kpIIWe+lc/qBOl3bYNDZDirQJKR5RHsAcl/6Sy9M6n7OwRHrMjDcDccNbSB28kwu
fQ54xBsFRa4nyehwl4NG/fMuOtJkOCzcyUt565JfntJpjwiqpvvyAnQNhZNXwXVyFZWqQf2NVz+w
+L1jPNsU/BSjPUauhijtRqXNtSWoXp6V+M5o5Lm26Q4rZY1MtHVzKlfc2S0nCMwBccf8iY6PVPL+
68wKXGtlsZYy5+GN0Xs0empGn5csxbpWF+1oWe19QN9mktqM5ej5v2jQGXxA3J4L69XhgS9KfgT3
h/Gj4rNAjwjMCcRL90N9RR9PNnIeO2+N2WEetQZLm1GtifZ0QZo+5/zrk5kCfNASG4R2PQaW7uzL
3i0HHd+3DFpQCp3zaxSODcBwu13u1wZ7JKOe+mNVngamhFRWc0yt0yBWIBG0ExJjkXybmDYHNvwx
NLJGTfGK72FSlPinOmO/vJtmFX95SgJVx/TQiE1Nojg1CxscPus+gY9/3qkKbd2jNA4p1tJ+YuYg
ZKpHfq70kPHVVSvaFF6OvLG+fVLCUrcIKFk1jwZzk1RtKXKddktPIJnCrxbRV5hyJejSjJmPnRpe
9IsgiAEzl71AdVIIrw4a9lO07aCgcPHNQdi3XnZYbf1ywgRpzyVD0jvP0P/u7c54lDZ6UKcLIYZ4
4Hri7M6jyDHrUjYGp3dpErfbuvlAiOzvAdCUtztuToIAXgLcAOQa7xXJbeVXGfYaMzovPRSXcbFv
0BU+cQgYTtK83CLAComS/wgPWvW9kPXBVlHMp/kDwzJFCzCgoQ5AE1p0o44ZfRZhQosXaYjDFZJG
zkqlMl0mgVBNrfy7koj/WeCffqIUxKSsHRaev0epZioGIK6uBMwwyFQTYxvW3SdzVZ14s0TRo1xa
x1BpBbAkv7DTKenl9h3oq/wbJH+NuwTO/W1S4xiG8EV0vGONXjaBYqTZvTkG1ZfUBAGyiUpgGe2+
ZZSbSAFoDAc+6fVBQBwUCT5mfo9JZa0O4VC1tY3YaQzGVevPpmCUmwFKPxXAHdcHPGQp1OkTsglD
fq/VRZa4fbZmTl2K0I8HJ1oZUgIfiJmpJVf6RNnlur/9PKli7Qr1AcODmVOIGSZ0YQws8bjytq4L
F1CLQJGwwxMIEX9tXJiC3Fnals9vFmti1GmvmyGx3Ih3KJBYbtOGPnZb+1VjSy5cEvxvi7hMQgVQ
Ti3BqunfufH8zwQUQB4nCWbVbwQYX+nLePDTWiULydK3j9Mx/9KDEvLP7WGrI5qagEBf0XQHvyYI
JaDiSFbfzsG+NvrcH/wtQR/faddgdkR/yorj+8BOYAW4+5C9vizwzohQ59PoJ0bdcgkMFA9gt394
c0kJ2WIPPeC51WwwKdlOC/SBTFYBBEVmNVSuwCb8OV7TqaH1ShqoVHX+40zkRPjb+19JEWoKXdw+
Im2lb7xOKyeS516WYmJmU68eZRGRyeZufjr5Z7C+fTAfy8Lz1VfhFKWZJCMllEk9jg4wZYMdcPUy
yFlRHLX+0bJhAyuV4cVNFcDrzhk8SBTsXTGh2nIvadIZmkvdG7w2VCAIRpCVF0Qrv6gIPVtfIu0J
Z5HA7ci7IqVrjd+shF8GN/T5NnbooEZOqi/u0Pd6jeFogN7u+er1EHGOMuRekKd7wxeKT7ramlis
vlnfCGPJHE1ESI8IV7L87v/W2PAz7TgN+MBT/IeKFPfpAL2tXamNYmYCFiKT1NOJfjB80tazZDnx
DQHvfyELKgfeBBYjJbckS5Rvyv+raHahxFd8R0spK+fG6bIIoLL/mvUoQjU12rWwi5otEcsNu5gN
m/50UJ6x0cjAkWsdGs6ifM/cBCpEkeTi+8ui7UgBVTmdTRpIwE8w1Qyf5sTk1ZUHIW1ga/3+McP4
qqOxaJ7Wr9WfzP+uyEgX0IrsYWUicbpO2Am2o8WLG4mI4vLW/DoO2WVASR5P9NlCryqoif/5m6gN
LrAF6Joj9T9mbOTmBfzOlcpckIL1jJj+Bjcl1Tfh3ODWt0omUMtIofjkgrozTI9ePEbK53ZRMXKy
1gZSda0/vZKFBGfB3O14F4RmDH//8JqbPJuLKubwMdcxEaUlc7i1TyMgfCBpa0OoLdZPiRMFN4d8
PrDWcEVBpeFhkvuk4SocGbJp4vPY0MlCCh6i971TqFUnvfn2eALJ9QMhA+z4cSDPg/kslXFQ1HSU
SxAISCWM7hVods5mOc3lMMqALims6m5gcuxf6Og11ZLFrgOFeBR0qr8gJOx54aqpyGsck/hiW2Kh
SaJhyfGLPA0DPLA4duAa1Dqdu6XwcHetFkVcpMTGQLbM2zWt14Ap2WbfECFgljh4TnDz9O+p+zay
nP8W1T5DDd+91ddlODAIdLIGESrAQ+aEB4jjtOlrp5YrFhGiHFuEAlBCKaMjFpUPFHxTFIJqWY17
KiJeyROfKU9zkpafk/pUTN6vpZgfI4+cQKz9ZUA3DGDqei+S/uHsbLyT9+A7ZnMHL6Uhhsn/fQL9
cZdLrep/HmHU7j9puv6N6NR62GvCHDHJL4HvYdO415JHWfKDk4qUeiWYzerhIXB5se60unkOYpKo
IVDa6He0e+KUdRgqiqLlwbPLN9rWetswRooZNzx5oMk1E0yBLPxA7oqEoGF5gxppB3VFeN7iBUoL
K0seeKR/CBeMa6nc7KHUDyjwyj6nKL8MB0CXbUnT94Oq/RYK3Kqtnw7vrKFxbly5ft9hBzVd7bXE
PjRBqHaEnzgJ/HSBHFppBzoCv0JYXhHKZaLBRItOLoV9DQSE2SgVZ4IZOJLTBoMz9dK5MVWZ2jh0
bG+QSVEpZ2QRVzF489+Cb8w2haxK5FeS6OPcoretYzxpN2dPuNnYaQz9YCbADC4MR73pkNEjZVsh
czaLiv1mucQfpBZQroGIDZ7V9t41FYceRUuMiQAmmJNoTb994x87aFHXS7eGda1V92U1s7R6Mp5B
pSU3pwvBK9wPj+l9kAzaCTFNgbumcDFp/INnHXxudOndqnlyeMamU1BZBFUpVEkRRmynDIFkMkum
oYbXcgLMVZKCAi1/aJDMBCcZfV+FpOMJYalKChbnM9DEUp0SNeTUA9sorB1onbVT2YGG7ghuYjUv
vWrRkHe8RmZkaVtIw47oWjjLGtoMRVNXq3Ob+m2QYbxQgHnWQqW0banfCFC0ccxqYGq8u9H5uJtr
S+YgCJ5KvaPojt6M0DR0oKZnnBHAQuGA1nAthSx4a19eWkkRgYWCpqTpI8xliYblVAXAjxudiymF
jJrSVCQzNMH2VRX1kyUw0ngBBf52jAFn5hwHqOulAF2iRNr6ftYMdwjkPKQWUpXDKNrVgFBBBV29
8Zr6bz28PlI6PYbEdMrJ8gbvOWd6yZ4rUlC+aAUE4PDDykzsbYM0GMewMbM/cP11bytD3qygh/hU
KB2zhDAIqK59ZRhE2OQa4wg7KrZTHooiFIJLRvyj4rBzCywsYAZ0RFHp895wDyEnBdwY+cYkrpk/
tnCAzcAQ6V2L5E/kM/+L6PZaROKTW2rQKSItgz23u8BA/LTWC+B9hyNPuGxr2EUiHNu4fxEjnH91
8QIg9PKtTSjEIDEPPHp3vk+n7w7sEN9LZ8OenRlmsEDlfPVn8N2/iheF3ohYsIetz4PloL40nYj4
vE0x/0SXb7TaXoELEL88ksP25nJjKx+i8c2lBWed3pfj1RxK98VV9a4/sNTOfsftpxBIlG0qG4sP
+DWrLKXCHAL2+7QfrW4LemNiOIp0G6K/W61MXZho+gVwU303ok8YdBAr5u4weFG6+AYMYIWLFZaO
SgOB8uyyMjUOI0n6uhaZczUwQ0h+xFG6Eg9fSWzbGks/bWL9vxw/UOCnBn0oeupqRIuhy/V9qkRd
qp7DMhaUTq4Prjca4fkBnZhOLdbsuEgJwot4hmPMs4a5Xnrft6NWlcu87jjgDM757uIM32SqnYYN
nbwV9ssNMbB4UZuM2DJsyKGZkc6XUaIjlVbyjkShdk+XwQByMSeQtwRCKgsOrG3DvdgFZKdbSWJG
KFua+QtUWVhPytOmyFid0KNk0Ai7JUJuWnZ9GH17u1j071pOT6e8tsX2EoCXu0veA6Nv/skrZGWG
FA+Mc4Oxk/UvRZ4ld3qq6ksG1Vx+Ct4EpNghvaG84a5OJpR8TAaPNUqSIyhDgDQJqytu92SVMtjg
vnRmX8fbLQIvuuQFpnNHbhXmC40/kcSNaJd4BVuvbwTzgPXj/UlcpiDqwAr33iyKQHp4O5XcgQH/
cgOobzOi+1Sl3OGgD17J10M3PTI0umW59r23MXs6uxFqLpmeJS3aqd2HcgXPcXEXpsV1CccA4yn5
NvbuD+8y/wkIBmxE+Zw2dY8116781nPTH4Ds58/ZrIZ7hIBmYmf6WTbKirjC0Uhfe8CUg9Yai3q1
2jnR9p446cFkci9FJrXOLu7g1KWqbIx3XSt/Vk2eqvXriXEQWj477f8WqDLI47il4eY9Illd7qxB
2OC/Gd/Qch+ygbdqdbqHaJx25rdI59KH9PpNG0vcVkhZysX1PCCUPdPePUPmbZSqp4RomrHr/uW0
U9JjVNO3qqh6GiNyK9WZFwoIqvPjlWalJV7+F3jFTPOhtkABuoOMKz9bIQ/GkIKwHf31t5rnq4qv
xsv9C4mh/qZrjhXqQLve9i4knXb9uJZExiIrDNFzHc6Lm99WiKaCngkFfaofyMdVz6MbVd9DjSg0
D0mY8Vzv124w16Zt3c2xz+doyewUT6jenKz7BJNbvTKwegBDsWxImtZKAg5NQazlYhTgEsDNzUWq
eY/SqPsGDpeHXRwoL2LXTJHy8TXtP52UBF5DDxCtLUePHkKKuMJqV1PMOYgAxPXB7kx+l0fM1oj+
32JKnGgZ+KOqutDOPZshGi304Sg1W9K8NGWfQnNmFGRAP9dX4nF+lPEbIM8WYo4IwH74jCWwaIev
SKpu5fQlCVybhtgp+i56rcjTU0GF9AsiWQXwy2P2jsqKltrQLm+ERSPPf6NbXpbwJU8IALzThmw3
MVwu/MTQn8B8PFiyy92EjtaNHSEa+fCDHBZ1Zq71H/qg31A3bFMJgZ0r/UYowVIJWYblyF/XhR5a
cazyeG5awDqdf3X4HYkkga8SCyFGqSa+A3dk13KTAcXGlBpBFIpYM01ZdrwJkcj02PE32Sn5gHNR
OHADNm2nr3A7WljTUkLy7lPtFRndo0mKkdYgH6QMEjHNOMNDoNUrzopEvbfnfTdkDSuC5OHg0MZ9
ZDDKFJ2fSSKPBPixQHbAtWhswbMykN5y6X/2L+4CG1oxv51/Sy4ud9xMFeZ0Tz/rk9IVEPgUn37R
lRapHwVERNuhIQ4iY16XnUDaYcJG7AqJdgbhyQj70wjqalk11Vs6buRvVMozGpGrfLnpvbyJOIkm
cA7GtXC+Y5lA9rKes92P8IN4olBHAr6BNrb436GqBCLR8Jy/lxgemPJX87Bhle08/OBigsaJrEKO
KEUNraeY9Gx6aBkbQ9pbrLblKgCMpv2nRAeMPCwLlqwwP6kTIx5kpVNjbXF0COUpjJxSIa4Maa79
/fK/8MUGZho8z4+63kl7Izhs34+Qokd0UfmJPeTuxRPMZyyb0JuztnPWoxOv90CewBkBvlSMcVdl
ij/dxwcmqGQJwsZ4uVmDPCXkxj6Z2NW9GvM1KGKQ/lQyUHLuEjG/l/0KNoJiLMt3Vbp8qpH5bK2/
v9omSCU7/tamGzNjCZebpBOh04x9vBFrClTDwkrQYqbtb6Opb7y2sEyp4TLFCu/uoRAJjka1ijM0
PmlhzQ38VO9HSHLGDk93nW7oFLQf37g2Tut6obrql03Wo9ciDBbzhq7dYHXilQFtNQD1mqFF7LJP
KDIBiMUUXGuYNJsnQn0R2XI3BeC7sHp2fsfH7/FlSgJUq3P15bfegQRAmXOHjWCfCcQNS7WOJ5cx
sSuHOUDBRid3hzMn+M40EHFl8nwZl+QOjk1Xv2Nz4mdaxZLVamvvKax6xSM0G+G/qnNg5279ZKeE
Jqqsio8sib6gE9mdO8AL1EAFXf/P8Afe7ArgL10j6hlf0Z98S/nGz9fNh6FoyU1QoROw+bxJsRwq
N0E7x9lCYEMyC8txWXENAMQNUsTl3opZEj8GZCo3WwfsgaIyxBDySQ1ip9C1SWlo4qzbPvqgwnyK
sPWuyVxKE4i9S3KH8JXNdCjIDoaxso0jV+/j0eB+NqoeyDEO4wb5LY6W8sL5sYG/lOWYRi7eXoQn
n8M18xQ3nWTLUiwn0zAW8MeKCv7EdmnU9pyIbGts+w6FNm9w1sVCN6+WTw19gtB0nVSMJ98+juOQ
fzkvfI/InxDuZ25hGNX7I+steHdAlQLcfRCmhqHju9G6DfUJqgEsqKRMxLBwALbLzqXH/vgxFXUw
NQc6877lNVOBpBQeXiXzbCk046XkJ8YK6QDMo+Fvw6ZUd33q+/dGOOTa4SWCMQ/+Zx7tTyO1/tip
4cXZC2KpO88WbeE/puV90/Fa1gcTLep7wdyOkxd5gR6zYb0gPD0bzvq/p783V4e7sfG2r+41guSS
gZHy6aQRhq8qq7eGtr//QK04zvnMXME9ub/qy9qjOrk5SDhKXHkIeSTobTLiJDZOUn4zupSXWlfM
1xioWPCkN4qNTLENcaxhysZ2mA3kkLh2SmcLz9fqK2Wc+/0ig4472vBhI2g4sTQCTOuXbYzfevF6
TQzYQlArbO7RPo4RFLlerK/jPBdRhlWWpAOOR6jSCfX46mPFoarH5SX80g7uT9F9I3GrSz2aUzVj
HydVk3HzHLBTCGAPRrZmRI3sMUIQc5BBuzXBXYce5gdJLLLl7VZgAtgtqLUAIoMOT3MLTF5qWZaE
65VUPbfhOHus8HI2nJbjziQH7RNYAXGCZoLIK8pFGs0VjMUeAfHZjTwnXwNpV5Anm9I0sQOxV2YZ
6OfHEVUlNcEBW9Vz7KLfCGH7k97iilmkgSYC2PD+Qu+n8ifdDiecvk6Rr11btQSf+ZpNm+LrQiLG
NITsWyu1IGSfvELd9Ys5AydiLRp8xPLSKsK75pXfemN4KgMPmIQrSnRXac7cDx/ZdjX38jI4iTiD
MgCBpHvPDnGTYGZlg/vPgf9h4ceYARrB4bXlwZT3K4x1iN6b9Ttx/2Ie0fl8TVTqwGnLUD6uYNDw
b1PYiYqaoVdzhFByapFmR4GQCO6Hq+qfBB49nocQRVYqA3X+769fFO0J//PYBiZKw9gC48JrQ/C2
A70XO2lwkuUKn1tDe3u241drN0XoOL5t8nFVJ5VizlFmUz0Sp33K18D/zJVNoE5DKSlpNT1/hrFp
nd0QI/FFhjaJq9xZeg2xqdX+zbMnVxMmlA/HrZM7vqfz8+fK1K8GNOM9+p3dwgw/dKVhzdUKatNP
U1YBaWadKIMxPtf8+XRWL6g7QLjmtTN3bIn5XK7WO7nlqjDFFyYkwdYL0hj7RwM6kL3nXJJ9sN83
2jj17n5t6WwnQo2WECPSDpRQP8zaKjTC9Pv+JfcKNNEZkxcVs8ZK4ouJNO3EI68CcHiaB86vCgWN
GRC6LA8q26ebyUpRiS3hZSJjjfsGHSthQJqT9eDLmA+qMv3epovHkGv6COHZ7qs0RChpr2SdB7vV
qKfoCn64GpW4CgNamsOcCqNxX1A/moIo5iFuyllV0AxT7WgUMnTuFXe85XLo8vv8CjrECIZ5cVle
gZPW0P5U98d2Kg9dxZe+f0ECxOhqyDPNg8IDKt2z/qx+zBJc9hJEPlym9eJRD8KWeB+mls6p+hgL
pZzyJuDx/Zvo6jxNzxgRQJRjsbPBiU/TY3FGIkPx9NnAyihG13VQMZIr1aCzwn5t9gil4zrUQuNj
yYtTsi4YzTAgB/mCe5cwvldbPe9FatbzCv1UUmSDGnyNFJBQCsWXENJ56uZ6nFvfZHgTIuRDi1du
3RjX0eDkyDtL7grl2mihXdX5IUZ3VZ3KSJJoMAPuXDWSlUn2HnNeQXEIIGqb3GGwXUcP8AVz2Rhj
on4CbIsnhnsJ6qozzPFNZkFpML1p5wijeDs1t09r3QCd2HKdwLSkPoNF43cVJi1ExKgPAyhvLY6o
HLiD2w+oAeO+ljIVMdijl4dl3KyhNDdnYQZiWuLCqoEMebxhvE9CS/iDzlKCL2LQ9VBxmyIF1S8V
S1W2Sop/FpyVCqqIEyLje/yBfz28y5Ryo/WWjvbW2TMjbWQ8EV0BFgjGZtKNcX+0+MTv3Wj99+oG
ppJa5dzVUF1ltK6gl0rWhAaWrwlrb6mtEWjpQovRPjsR3EfMuFWOj4qU+lUYHZe3uDEgibZICqgS
lf1hUbcOl2/6+1lB6WZK/Ly4qTeCm3JW6ijZUZZX/oLhU4+CtXGxTruDiOmnwjUDpmeTzm9WMEmw
LsJE15DwZeRlfR0zMud+poQXgkNGWi+THuQr8u4ZDrn9/YnWKdbr47A+P0nJXhEfy36A+mLHUYoi
PfnjXf298MUwGAH2odPqFiXmNSYWdUbfPWLMcEGm1C7tCgJT0a1UDq/v2Ha0KCk/+eCYs+4DODJ9
ZYEjVEGJ6WnvYuGOUaqwvZ6lWXJYkgo15mOQfoNavB9X+viPkF2UwpU5DLhHINzrizkRS0MjcAxE
zeRXQoHXw8Iyk6FiSUi4N+yk82zhhzp612fiPaxa3yHNbk5Tz944TBSYFYuMZqrZq4Q5OYgNmAME
ldvt5rlzsoiI3B171M9kDywIorzuZZXaequib3j+efBQJRJrgEX3tzvjV9AJ+Pe3hiZk5kQS7Mgg
p0FL9FFAvAYJ30XAlPHQkIBhEmP6ng257MiFzuaEM3C7LduLFUp2CZTeUHni9pxgjmoEFixzkege
SuXLYNbqo0SRjf/ZLfDhlSpwgbotow0mQahVA5RyuNmDMr9AXAmkeX7u+8d7Bz4XMmAKyDp3PkbU
V67mihxAC7lVcmblpoDVo/5FB5zK5Wx/7qHWxw5qhJmBV5hqfBzJVxhhRCHs3/xLPf1Fge80T88N
6TsT++FQDY9YHL7IwzLSwcxcRA/vZRBH3EFSXI6bY+oBYEWj6OKezE9FKtIoHDZz2dkZtXiNQsSW
onmwpAr2cyX4mnyrJwUbkBbo/UxR08uhLxMDXoj+Xp73m3FG+5h/rQMY4RDy22WLlyWMoBHoDvLg
/pPUGYoK8OvKH9ElFyq7+RtCCY1roeaRl1ofU5hhzq7Q3XApL23FFnrApG4jR6fhfr8m0UUsf3Of
MKss72Pp8SrrIQ2adQx28gm+b0merdq2UU9XVMjGRGfqU6VCgP4D5Gi8pNYQ7QL0tqFcFB8JSZMu
oBNphartov2n4ghDD5J/M9ZR0o2UckiA3t9uc7B9zdyUqneni0LL0rqljfJL47OlvAHsTcDWtpNd
UlgJ7LtxBhd/JBbD829u/S7Ho3EqZE9vnttqHtZhTwsYoMHhqAwmh1KjWYnHb3KUsEPcPzZjzTc0
+0mHid3qsq8iPnXGYdjXNS6DV2QKeDKcFxnPVW2qGBYME4TEj+c+ZF2YisON+OpzM2nOoPc8aDgu
HLTcNfSfg++NLdrxF2QitW+61cTQYwyMau26ibGkSJ9MEQnjKvibPp+Wjc+pZnqH1HqQJkdjscGs
HYLsTTFBLHzfiw3OuRC0mH+3uX5sSxTQWgxLl7SdZaO8tnwY8C1tBmFXDarLv7LbFoA/Tt0UfgcY
DKlsuYy2sUDBmM3wDbFQiyru91hL8jekIT84cpptfI90cZT4h39bzUVUntWVRsrg/vmK1FRniVh3
2EmRVADZuH0dmG+7isQqK/YGcmnnWVgKcDSt67cxFdhtBWaqoiOkm9pHDMMkijldraDFVvAfCmZo
3lPu5bRlS0+CUuQQh0/4QteIos6O4q11awAsEmWAEx/3KJnUvPZLzWQap6guDgqrZmb+rFC2ZSoP
KKEkPLCe2TIc49MJ0YTyVy5M+HycAqdGvI3jvOLC7BX6kvE2MScs2MYhzlWLItcPUNT+464lverh
hw+4qRVDkITHRWU0hsmcP2F5zkowUvMpTAnz6ZXu7FeeYT3nCUwg5XPrgrQMCPTjL95Quq6XPcY7
hemWUif/AkS6nEJ2CgP+eu0KvTFQlLNSAoOkwT8g2QdVVO0KlFFz2S+L35/vtfILHFAdabwg0/bx
O6W7ngmaNKxfYYcyZZ1TdALXzh3RbHG+oloQR4gpn/kZqpNDmZ8ZrVgpEaQAoKHLgi5GqmSDq/AX
rfFB+nr28CeHyPxJA4vyHJgLukMQ2YmRzzzPSfLld7t84cLlftq8FzB/1GxxQ9uihBvqfCOhi13h
6i20Zwyyp7vDut1PrHF6Uv49MrWW1CdGEKUOhSapIIswDNUl97/ZE2eg6WFfPJ/yrPDKZ+DW6E1q
5fLsqOJW1/8GmWxa/a/mQJ6IJvCKPGRkBlwYDkPWIQL9N6iBRdrQGupTgmIOb4L0AIQSEXyT4+Bc
Tjf45idozhKg9N3B6oDGGYt7d9iGI1sjsyweh78aSP75tBDE9rElPQHpYCyhsKEnr/Y/LCR7p96N
ZFpniH3nucariIkUOfjy32WldR+NwyfwR0XuM7Lx4xyBsBraelXOpmdoojs3Jc67Jkr8rhSSsRF0
x2sHaI0XbGoUiOX5ppEK2g7DMTyrzPa8SdZI3gejM2vtoYpj+1yzFQ4d1raZUeHSyWX334deWcfZ
/C6CcHzyQt4cerlex4ykftHiGL9kbBS4k/v4Ei700vNwd0NvaHnFLAstHnPcpcbnjoi4Q/MzCnB2
kSeP3Xq4HeJ5ematOQVwIqR3W+mBKGwaYCKGI0twnEVdOyk24oSiRbBk205qTI3ikqRRLYa7/GHn
m+FL72ACOHOqfEsKck7zaKTAwQLhEE3wXe9OUdUlP4nx8uyb0vB5PMN0tDco+gVbOpePQ+IZnB9a
8XjyFFVipYH0Om7df8WFyDNfTll2Yeq5uOj3VVt6jsQmOoWy4H2l0UcUaWxuidMuO26rmw73BG08
VECUelGf9S2yCOu1w6RKcKwZgMSSU5ooP3ydAZn1/2DQb04nH1XJcp0P5e2uWSKUSEBxVYJGxGFX
LgdvzDFJrzgRe/BpAAl+jsm4Cqn9HfjofdJftI4vwrGkr+M694YeOcjZYAac/Av+QI6LOTpYtMrf
E5GCFxVQFUgTCvXv0VRMQ0AciuZvIOTAiwuMnL0XUCMaP7e6A5dKoflNmdgrjNS+nyhuw0QxFN+g
Z9AQ+OuYkUVKUP3bZaNTMlGzXxaTksYAsKfl+Ft3t96P6t/tXdrgkasuqcmhRt9O6BNDdxk88/fG
AHesc6XweTYfe/wYDZfRWtpOoXlSvWV87Y9NDWwPsmq7dXWYWi0B+3czHoQxyNTDnoxGd0OwVieB
7lo+DGO9S7x81ZHYKLQItTULHMPYAraob2ZSKl7ftYV3NranwkZuY2dpLt/0pZu1dLfxw+0O9o2p
kEBV9t+tgMV4QL09FBa1Rw63Hp4VaLmgtWzf3kmtkup6f2uhQQUCwVWfbcn/jddWXzetc9W+JSwl
64Sd00q0RE0RS0uG7Qri9EdslzsUVB9ESjklcgc/uLkek5VjrboG7ntUwAJG4B10iFYEsSD/Y4Il
zv+4jqI2MggKOEnGgZr7++tSEt4ltTM6OuNTevAo9F4EJ1VSybUaP2SXG5QS0dM8sWzDYes20BP1
+2dNV8iVDXNMaEUznIEJKXmH/8TIuHylmDt2T39FwnpwrlMFME9NIWgvsScmsyOgI/DYF9C/I8rY
qf7viqbM/tRMoxnCGj/CEAe6HwQq78ssS0bZJTh3RxYNAUBp+Kvr+zffIcSNrqgqP1YaY7CuvDUU
uExrhP7uqc+Egzjdh77mU3ZNex49QCchWjAzfOFIjeJFR+R1Fd2rdVkx8nxY0UUOTCnvxVrSs8UG
sqBT5CA7Ddn1UYSvqmlaHFdr62uDl4rchyfU+2ydgbvBf2DPN6cpfKi6hL6Ch0MPCL9BCZZZosYu
4ahCtjguk0UyGw241e56ze+miC0gDmQkmXZzGUpSfSVvK6Z/JKzuj3ccmnRcU09GpvIQ0d7DQF0S
UMnklJmQgx5Oymo55qt9LPvD3/oJ7ApeanaLAQ5Nb4ZGYLy8FNY1MWD8ZG+Xaw4f5zaeMCGQoPC1
tavlRQEc3U1OjNVK5BJv7si/ByT4xh9bSRps/YNK0wIHWVFDX1vIL+rUbs8OFi0rH8oPUrH/T2Kd
M+uBEa1kU4Qg0OTfFJYOYWH5J0ZUvFS75unP3Ch/lNgUD/wctMaN48NatMjOU6hRHRI5Rn71npDJ
qulBtzKKklCm5EEAFATeANr6td6saIRXZ1rFI4tkuasInQr8LkAo3lRTcsmgpOzzCC6zWJIPpWii
NYQQFoY47pKR1gRb4wxbVJwCB+pnV3pklGfuZSKR4SNWO+Zpil0mDDUbokx7fNRtriwig8PBRUTT
pCdA/S7r8HzVwyfzQKPNYWCN5WQxLvxrQzv1Vu2bl+F3Fq14l0NEtEHMU5xk0P84boe2HZ/Rr/2f
j1O7mVCXL8KUOqguY4T16uo9/ak292Rp5KLLg2B03w2QLn7oXQAXCkB/ijCL0sgbUp+6AJZmjwEQ
Ma2DnRzdp3ROrsKJA2CgP8RcVgn+SQMeuNN4WKPm51bEVzy+SU6OBYkUKtg0oxJJYAk15gP55A7L
u+s+vsC96kwIJnqpG8MlphoqxCbpJ6G+FU2x5/nkEwDpRuAXKPtjTKWK8p7D5hNGHXEsHKuCgoY7
noIzuhi4/HCRPuWvO5OWbPaZ3ARaZi9CNAAnr3zOIj1U+8PKdj/SX3MVzTd4HZdS+ZFEOhjhyq8p
QKBqd+iSDd/2eO75TJfBneO/QFy3RxX1Yvhmwn9TXVMyG8+QlcLhzVpAEWITnoH3l8KzsUNbBDLk
G/cSW9xbOy1hM0/4OXjwxWRMydZuG/Pf45Iga5N8DcS1c1VswigKzrlDQdoswSp01i3yf2YARSUs
+3yDtc76q4k4v9YsYfhTkpzY/i2Zd3CgGuzRH7EF4S1dC+FOC+tHxq+jnLgYNkidGvrN7+3d7WSJ
CdoCVPqFpkBjv9pMqWRZiMJo0genEfEv+orojwAZVqVQ/NZ0/cpKgf/hayI9mWBzOXRi/R1bKiA3
SgbtiIn5O9UX5Sp79dblHh9JxHBg4DiUe6uBZuy2U04Hxo17c9RDYzjdRMrOwT4N0OHrni0y2FL9
VTPHV28o14FtVR1Fnhbgfpl/2YdLBHQE+Uv91pP7AIZQvGfq0G6wWZeLEFpDktOHgOObmsr5M66s
RcovpBbtB3wKFJoOLr2XnK8YcvEsrNLP5pTwsNJM/vbGXQdplXoPmIivpn85uGNZ7dmeSAuchehB
dTT9QTo6dDZR3iuBEE4EVu2UDdBPLJ9xGdFJAN/FgBYZaoaZPlqAGOWLujRGjQs7/XedkvE3BXwV
9ve/9yx+GEr6FSfNFHCqEw71j2+eJXEw1JBgcdCI1l8N9jeNeAjp1iCS2bQfzbf2QYnjKkHS4zyw
THpxZTlxHvid5EhQQEFF084e+Trd9x6+/5CRXmARSNkyrGNPVqqqmNlpucpYbJ0LhRH14rF8FHE9
e4UDE6WN8jqIUA6Ym5f7j5AJLcTMpLYKyDV9yHGyGrEYq25qDx2H9dbv9MtvFh2lVikDbdeVy2Hk
iCgF+T1xbMx3Zb0bmhC2FAiILCR7sYEgf8YAAdzCLB5WSAvglNBvDk/ii4nT6RvzFzDTSnYgvvPZ
6BgoQVIbd4gijUgu65AUUqKnQqtoLw55ZH+0jSgdXGdiTazKvJ4WgLGOY3PKa+5A5++W8HW8hK7I
TuA65phz4ze3FeweV1952S5vZBlKNmuARqA3Qi1JihuN7U1QXUHFEALreyx9wR6xFcBP4pdhSQ6f
p6QLt6whfgL4wg5urN0gvlv7co91stKLJB0fVxSXOV+Qz0R8A0DCrUSquyxW0zFfzCWkAZn2YDIo
YzZs9fbGSzDJOhEJoX4eqGGIFDF4ujyKv8xNXHevbFvameLx/xxU3VyVl8n52AETUwH2jpeebq+w
Zes7+RBMGLObbNTn3iCxpf3RkAFQHmNTX6y0AC1lpZMOLOnq2vmIFDEv0pMAQ/4LCV3REMATIURO
/OKLpGX39FhgQZI0mZD4mGg+CoK/lfU0kvuN3xWmoVAZccVsHxig/5NMvn9xraqlygRIHiLdCX9L
rKr29EOm1xjijCInkl+QbjkCsSKBZldQ7dcOCjm43E0IpF4wJX7ieBukjNF/g6OLs7oQLCM0aLFF
MCZeyGLdecE/xLJfzKUzxIsfQsX8SGtWvA43Q1IkibwfQsLLUeJqRI3bffQtUPcxuVruaTwo0fkD
ZH1zzhteoQE6A9EFAXptKfFMWKWiMLj71oWtCMruUoWmuKTpyLz9mDfg9FAqnBvHlQU7O9ayCFkH
15dp4sfMuHHgO7kLv5wB1eBYzvqMC1WmN+pzNz8hGbABYHxciTm5uHw3A4b41HLnZvej2FKCLaXt
rENLXbNDqOYFET8zjfvLP8erI3ihrKPtdoYFv65dgElb2BENVR3WMYusjP67xO/10ZblnoWjGAaI
fvG1ar0QI+g8EWrJ5JNPTp4ZEE9+C99VryjcvmHYCPPtMXa3GYZhrW0h7FnDzniTvygA35/cKxwQ
LobknxgeUl33CQrKX9/pW5BwzHOASDmxIuExIJ9XZtB5yrkThgqf4rhn3aa3I7ydZVaFAMvsVaw9
vaKkAIU/F3aMmQQ+RCwrbJKOMMlXsOgv6BI/Z9tkEaZFxJUpu8E8E0/YAxHcQ6iWS+LKsQ67Dtqh
/4XgwsA6fpLfIwwnxXpPIB+/oIUv9EMgub7BFvr2951u8o3Fk5psKX6cI5xntqFPm6EzmpsQLYdt
I6UG5xOG+ZEFkE+LjxUlwdDUF/U6g04B8eti4qBtjTsEyymgn50pr6IpoEehFqbTm1NzdrX3slma
gDGukumAnq0vj6qXia/tulOyz9gveWQ5voK++J9cvmIGce6zykGoh/hBNjFteEtM4zz0JkLfHntO
05dJGdOTn8YVWuciiLEYdELMAekGil4bC/sUApc1LsMng1i2Po7gCQyao+HUcg6MCXD9rrrspCTb
nWYmVMq7zTqgaQobKnHWML+2pr5RFSUQPtVjr2gu5XUGIwtLeRp/RE1tc37P8GVUcDXh+nhAdIvK
zAXPhbVPKYk5oslbA9aykH/LEUH7i95XinHjKRYhGlN5IghD2gb4PGG4/Yr4F/5s+OxiLVpShBa3
5kRcJs1irhRrIFOWIEVclowCSvooTRMpBPl42chlGtLFcarsHz0vet8sruSx/Mn41HLzaCDBEPW9
cULaM4x2U4rOBQ2AHEM5eRH3e4w/gsxWOljCUsdLtPS0MvcSRlHWxE9ZnUJGtW0RsPUmPn31yAWF
YXx6ykvibTuj38jUTgEtLZbYbgjmBrZ0TDldEeIfuVvktLixTwZPPbt8PW6Q/I9LG8X/ED+rO+Mc
ThyFslphyjQnKP6QcqUU/ghaMKGTAhMWlODhAD2Lkpfg1JUwCXVGxR7A6dmYwKrRtQZNYdoEcSRx
Ky4xFPlrl0U9md87VCyawP6167f4UtS05a8FalmvYHN4m7f4V92JMIHI3BCcuVcubM5m4GqZNM5G
BDij8lHqEnOVWMNmrG35wMb5pYG4z1ocDh7Z0S2H7S0VfBGg09dJMasIPY/E5oUDMZFgPAsYnCqB
lK6tAxaGHvHXHVp9NfUePNd/wCLHPX102T73XvdLIVBJWJXecveCO/wpePThgh9wg62Uoz5EqVAm
Id/Vb1bJbcyy1G3i8CB0pvxsuLcnlv4DsIIFGC9aKEOeis06TfXc5DrtnAIW1JTWLn05KbXdor3b
ENOl1NoR+GbDOXB/6bC31A65msVASG7tAx4AMBOr8W0KKfCwb+rfBONBIfo8VUoq0dB65lA/Hzyt
h9R2yn+BCrQdeqrRAU69TPCvINga7MiWzU9J4crxOcS+DlSSeVXhlNIdl0hrQO1n7QiQToyH+kY0
45Y/uPlSQx9RCklr+qMnIQZ0KVi4s1h1bEWejgKORAnRrZqBdYPJBBpb+fxJ0ruGzURJdYDwjsvh
kyJtDsoURitYqXZESF+sZ+FHd5HJ9zNa1wFzaYAupDKgsIA+2ZXd1TqYUM2DXl/D6RyaBtoNKBNr
J3IXPpE3J1aQRUbLpH4hl0QdSEwDWc/M4tbfHEo5/KZCPCzqTtEwgF/vf+W96tM+F7Ep1DjDipJ8
t/6BmL7ppydtnDjjyPBeFdl9baFww+48jnCbGOX5tEe/YbN8h6doXvlSV/LugH4yG1Lxmpl09w5C
jiERx2KWUvYNIM56Mr40rAwM7nsHAtfC7/ToyEQc8TAqE48NOdAh5zdvUY5ijRF7afRc+1BqQfzI
u2oUE4eV1Qkua0QqLmIZNuESuMTtL55zYUrREQGipLzx35PxVnnmR3N9qUVbnfWVMUP64L9h1Qvp
eL/fcAFNFlgZrFyGwibdISuDOnTmkFKvR8w/7+zUDtwcNLlnYmi2pGykigSqlu7lms4wZTegi4/J
xEvsaPffHM7wykrtAbUcsLg6ZJP5lhxu+dx2XOejJR486YF1PR9biDabuJpdNktbEroJVzhPoyFd
Nu5PEM68+Px2MLsyeYeyVAYKQE/BHtNhvWYV5EQug4BqB7tDV/i14nE+d1qGtE8lk1ma3YmeCoAW
9NOdAZbfYH4re9pXcBdogWrisuyBod31zMvF0LPPB13sQSGAOeN5XU+7uHeeQQ3MXYv0NYJ8llxh
c+HSDX3PikdonEIReybCTP7kihjUSOhLyLmPYd0FMzJX5PEpEQmPepUF1ythMa5AUAVTlezhOv7t
nfGBw8uXHQHFbjcmmfM2PRmNM3Tl89Liz0+BF2hCS6rcxmi3V8gSzGoNppXzZ1PhTgsJKU0qE7eX
qZRXShHR+aVoVYLgbHozC5HQvzKd5fIyxxMg7t/OtvlpMnczNU3N4zc5BzgyDeE9sAArjbTzYbhf
8jce5hMZD7WZTNkGxfD65qz4kvY1jg8Y1DQue/Ws1/Fq/No6GrDtzmS57fR/NV1uPbrtwGpcA/uY
KxxoCh3TEHOF+tfE/BNdhQntMuWj++aFtAjeIFha41cmtRYLNNk05M4O8R/vUteSlK94mNTwm/8P
gWLA1pP8Gdz4nAwmJBYoecFIN1eFyZYBjfyPF2rPAZjQWgV6ZTueJycJPraJJYb6JPtKqtw/gDKT
35JBMHs8aXf7Kl8TT1qlRaDTE7Lzw5G5VY8KAOX1412H1gBueQesmdlZ/3saLG8sKkXWC0wbJqaa
anloNSD57vLtivZz14F5Cg2nE4xFbbzkenWencG7jd1LyRaRCJe1ust2Em/W090TnhIGpW8Ur6RR
s/aDCWJ9HlixoUj6lVe502y4MIT9YSVnYbADZHm5KanTp+dV3clPrkGAlyFMZQBTzBWVyUpuxtRD
sVL2E6H25iCubaUSiHUN7UI6YdCKjE5CGWv4ceN04j8qbtEyAkKnRIbklmsLF3tNxMq7ucF94rVk
nAvLqAuRK7HxNSQmfnDd8bENwSdxSE34hAfqPbhI8xLnhJB8GnaFL/u2uBVlr6nvuLAVi0yuZ4bM
Pb1Xy3i9H5DscFuKPk5qsB+aYx/e6/LCGU9oog9cdpsxFoDfGOS3ZuF1yNZTh28kYBcMimIemW3A
accQGc+WHuj5uXnCMbaZLS/wUCeu9xq6nJKYa4jvloGV8qKtK0AADd1AN1OxQgUXi1vnaRzUTXCl
IXRYEQ/SSCUVglZXnDrY5P+DubcW1Ic/uzn1cR7YcMClvg3wCKld4D+CmtT1NT85C7e4asIx8+4G
XI6AJf1tQdmPVKjO6l42lVzJi6VmGhi8cpDdZq71IIjDO3u6t8roE8bhPU4zkWvXxByF2miYdHW/
4pygtUncO7ndwCrQyMjwFAA0TJsdgbnGrOYjQ5jOrHaVSmKPkdS8EGsxTAxGnB4cJdjnRvvUr2bo
d+bl7ITi2rvIcQS5J1zqI50vqzzNPqoeOW7bbtle9uUq03kZTzQSWf69oxOIySkhih5EJPbezpW+
kDA2epJu/kUbGmiI8l+DzbflRvy4O/KNN+SSoJFSg/VpACe8O/OrZfA7KU1X5uFp7WkKwvGqtb7a
5eEb1EBatuluPvd88MUA+OCGUGEBMzj4Y95sU9J4wYPCT1RJ54XUth/sbMtGJFJhmB6IoK4Hc0qa
xBiiDufMpaXUPnXCwWF8kxG1eJWVe/t4rcEYrXqnJp6CQpP7kjbIOQXpZVe6vsCAHlkZehX3QMUy
zk94vlfm0dM+0H5cd6PytCHffXRK/g+gcxiGHLrQoRvLovsr5oyClYphPLAWfrcQfmutMWJWt6fN
oUbBVQIGlWVmpmTcw8V3yEp+6VtJhTMC8aNTHMKgVZdghCwvksmZhRMte7ekejZ0bmTskgI5/vVr
7wdcXtYLWkGyAAHtZeaUpEXMewQ3Zk+ISz/TgEIzLRo31lH4vYjaP5mSpHq1V83y72cb6D/HgXEy
M4SoGwA9GFOW76W27GcQS+w21hHPi64Cr11GCK2IBVjV8zgAWdxQFweH8mYciP1VE0kTQ/7hCp3O
Ohvl8YN7pYJ9zPEyfV3fSP0kM3evqFq8yInGgMEAd3Q/vKTN0LbcIPg8aakBWlnGGxjOd0ePab3n
EHbAbOyhF0N342BLs5AtnmhaQ/UUdATjK+iHSnD1Lq0gRZqM/EzwfLptn6/2r1AGtfV4Lq0tY6mb
lLNAUD445DiGEeIsSkVuRccoi8IBrvlLJY8cB41iuUkHXRtiji9WXZiLkCqgpPDh6mdlhoFVcg4d
K7w6E6dg0ODiX8Sje6nJmLDQ7TEemlox5kOkuD0evB9dVivmpJEhifRQ+etNerh9uMoyp83tz2O/
MQKNZYk0a1D8aRIaKKP2aMMH7J7wPMAbARJ6ulNwwV4DUn4QmMUANnbq6eacWEVMPIpA1UR3bm+C
2BJWIMbdqmIPmWK8C/T9iwJ8ALomXuy865UciXbn7HATu7vZQGojd7DKJ7OIa+jqN9Q+Bn9gwtrc
GrVTVWu/myrFQ/omEInTddKOhpuXdfNZMFlVZopA7Dc8CCGNng1RmLUOeZFDb5kxZFAqXGlntP79
72c9gePfCbZnOdCIVzNjWoAFxXqeaBum/KFgd5jyznndw6BfeLO6fqdnxL8scCc9RH1s8CcgKnQg
Bt7QUpkwSKa1RCTGGSzA/wCcg8evlAU+xGkCVYWEbDoNjYYTLDW3MTjTOI32stVs588dIos5GZvx
sZzW8k2NKzRFRwNW5+4iwrU3//W0Uz0F1znvp0uk4ndzte85UVYWSXl3+ye/bBhGO6L2AyQzVFY8
FgGzUBUuuQ15mTKciVgRmQbKxqaLy5QDgSz8tnTcfkUDqTtpmoP6qaH+kUkU+0h600VIPlytUDuw
Wud8GcxnzdyhOATh2JyvaABHVswpC18DTJFHyM39emonO1YH0ivq5yOOQw8vFmuiLxoysfklilpo
fcZjXVvbmLxe6wGtn7o0xupilghzA0rt5Q1pt+kaYSeb6alBxyrW+JNGii/JoVVK34gzQemg3RQp
7nmBMsmupOeKofTG4+dY6UrF4MTV5lgENc9kXXHB1oqLZtzHw7vpAvgDSAaIg1zzTBY2B8FDVmz1
DqmzR8vj7xl2Xe8CNI8FaZtqwVHw84zT4gNAU1mo8F3o3St92yH4lswqAHm4Kf+SzwMwLV0kw8GP
BUp1pT53FuU1eUdMjw+Uhvj25VA+wqYqetU3Y4nQJFn30tYU2V4/UeqfKdtMF4E0pMHoE0ye2jCM
HU5i7cwAuZhkKvrjiR+HeBusE59xrnFIMmNSt5CNZHWVeiLdHpXgaXaxYQ2i7UPT0YM5iGkynt7a
wrrs8eaHB9iDDmUOkT2UQzpACR41K/HE842yCXyBcOABSXjvt+ArZ9r0ygGmz66JnT9CyGdxxBRc
gcADM9OJqPTC5/Pay57dq5YGlpMm+pg8jbZEQVNhs4hephxj8UkPALE4RIAiTSyt/Zx34/3IHWsm
ZIHpWszya/GNDZiEE86Ba7FPxoh0ciSSvxlZPLpVAZJ/I7VW4+i2b4E6jBoWGPRZEege3hx8oVyF
LRJaNcBUyACcDhpakOXgowxGeW83xTwp62ohmIwfdbqx8oUHFr4v2plbMyCpZ1qSMClcFHKKrPAO
xFJa85R8seBCc38NOnIXRGAbuZ25iq04LSxs1SAth48TkUaLjVDzphlk+LfiIlcdJmZtgxhSWMxV
qWxUsLdGUmHsbsO8dZBPlnFFASSfnqS/kkbl3T60jqWWXISpWVtGLOQPNrwiPFrf/33UASS1FwTQ
TnQk4X/k8sGJyeWq6yqBeRSnc10mNbKHlGoIzEJIWxTzc0f/YrpXsVC+DPISxn3LUor+6Fpaa6yO
MS3BywNDJyNk/PXQnS8w3bDfCiE038LZ0VFcbW5J5HVOT98Jsh5pq9+ZFEXahXS7ntAhf0NqabOu
sKyhyIvUTco1beL2WOAhli5zofiNQwChnfQy3QToz9A9YiVkIqgEd2aAXZydQ9vJS5e9jBEwoV6P
9Ke7W3987jvzBbxrTL6GO8v1kt0ToUngGMiuw2zgqpeSXK1L3DTUZfj9WtT5Q5g7NYPfsSY9R3Z+
TZZhcNcy1NA+Yh6VAElNbG6mjCUt8peTetTI9EHDIXNNHJiJyiMeDPDYbzImYaPrav+2tJNLMM5i
QMsdx5OQH0XPtg7t3PgNhA/hbtTO+FcoOnHbShrklWCyjzObnkCzPHI8BnKOEO/e5mupVfPARgov
b/n5rb3LuVPPltCRHtLPdgAhpzSNfutxL2s0/9X8lvuO/AR4+ehncxyV5gmNNBMXflnu9RWpo/fu
g7I+j6D8rg1uS/CrOsy8Y0Ha8U4Aa0GDXd9X3G9dHyKz2AikR1U2MNfGDCuaBABgxBTuVvfvYKow
OUNJ7fyB4J6KjtgN4799U1hV8MNObBvW1PA2nnuOgvDS7AtgfkpbQzpRWy3nm8hStZTuR//DaGwL
kvXXDEensI79DoUco99HYwkDuFEqAtRAq2uAjxIVabw+42OZ4gWSq9jYgB1fH+j+eC1rkL4qr8HR
V5E0Q6bgawaZk7chDj9XdL5ZBUHNaQevnHaEDDpaQdsV7GV9HxARee07SpppD3rP+586JdRlXGNS
O9qkNZkCyXzUoWpLe5+JzZbWHPm96DUAxct7lp1SO4KGfQ5o40pWtgLAF2sDANFeASYGgGLfO3+M
HyfF5zlHy3bfHSOpIhJ2gKKgmG1sXgCteWJOvskULKa3PnrJR7xwjMX2gm5JfuASEjVea2twaeKX
FPCSR/EKu6LU5W51f0qozzXE5ObX0Inl1aVRh4ZvzMXCGUlDIVfSHSizHdB1cpk5c34SL1E71EqE
P1QQlsTZ/bbekfS9EOIl8ZHs7Zb+bpRIqbh2c/Lbnw+kfjOCXVQjgi+ZFUTax7pmAImTm1of7GR8
L8wr7APduCqaHVeDBHmS/hpCMKmAGEhMrxHy7mey9HTn2B/GMxhCNVJErOW7SC5VTSb9XUjlehXz
6RxXkbIA553nN+DEbflSPaxAZx4/ZWHJvfUB85IY53r6WWCmmufEqxZcU/63gqMlNSYarvy0Q8kK
ureEkY7ctnkhn3yOXUypkRejfOM6hafkxpTCFUK/waHyy6zY0E8eOc/R4zjL63Re37EY4u/6KH4L
jyPB+iV2WJzYyVKKEoS3npDrmLQPWTQVx2TAWtwG9lbcLxVNIJCkXwY3Ra/edZN9UmSvi9omTSoo
FZQRnw2W82gg4BO0hAInwqGNGfQUaGhzjSHnAgG8mk/eZnP4NkXEY8aptOuNqQGFhphNGDqfJ+xw
At7BSttuOkulGCaGNIJveLfkaW56zijV9WsjJlJzE0Mp8/5ipfKGJtNVGgOTZdfkO4ylcRpCqIXV
3zkpYgNXFxmrZC/N6suQzhCdvvkpLgNUwgiO2EKyhlX0i3f6jgMSEs+uHgmS90ny/LDP0PTz/fXA
O51unixARYKMFpfHTbma+28WSNFx2ZDd6Z7fIQnBdPxDD5ewSPDMYQOJGSXZRy9n8ZlMBRqq09Qd
R4PuHh5unpUCq17Utl/CTCvEOv+ONKXiPNWWU6YJoSWN/cjw6ucui/n+eut3nbtW7ItKy4KO6eNh
Si6Ey+eyRsk8a8PmcZOq0b2oEZdtQKSipIV5exp4N7wUNUsCLpjKukko5PmlrXZMQtD8xA++CNNo
LQobiLtZzYTDYY8AohE8qRrrDe3WbyE8b0DF7etquuKewGNYlF6LI790G/N7gN3NOPZSED+FjOP4
P+GkCYkri2kbzLJ5okpBmCDzk9S63xtDvaDuA2iwN7JQ7MUCos5TmSoVbpthFfJ/U82r/eVCPQON
d+OpXuAKsr71DUb6XkoEOOwakzg3fslfyY5qPS6dQg+c89vFYpwUESZzBWzOLas3dH2kQbPUWGZS
nS0napvkZy8RccMeKDGqWCwckUHrrGEZ3VdZ7vMSzbi2uiS+3zj00UbGVt7U1KTULFamXNs9uAJf
sUFhigATXb8nesSZkNIxywkWKzu5uDiegjAv6FKF5HLzfyB3dFHt9gNk93UUrA3njEa61kIj3eTQ
5UUufJv+6BSC022M+7gBy8F37jeZGYoIE+ksNf8RazwzG62MzQmrusi7e2ej5PZV4LGxlPGmhm2K
CH5Nf1mXeWMpGg+OQMbwe6t5Kz4yWbfsRG9U96aMhiD6PH2SR25M6xV5Zj4qsi/qWCYEhbvvA592
V1hSGsVfrul5cAbyH7yy++RzZmdGmz838udghiLZY3V0q80t/liv8jwxuhZq72R6A62nBuQHmfUZ
rNsNXavi/OENQi2OIOhexysQ9eccEQfnkl+33zsueyZSsKdN/vkE1ptwuEFK61/lUDZaZVGwZa1B
gyo5oZHHySsDFrQzWZ4jKtlUZS5epcaKwJQx8QPa0NM7DExqNL4lZcHl31osiTI3y8cA2pVplPMf
xF+6oaQA0kulr+eZzOJdjCNpYEMeBqvNAsCRnK9SvulYRFEZdR92T9uxe7YF6tu1XBSRrQvwYqSZ
xunP1s79RfYRRWpdvU7aAFeoVIDIXtNOp0H1Q1OibCMKBI/qnQ/lgUUlZo/g7Mv7btlXgo6iynyH
hqoUcHBriJxNmOPmtOLKPO1MLnb/m8LVqOdDWwxqMrBiHMcUJLVhtQ10PN5511uFYGWnBF9W+huD
RaUJjM8wWZ2GtfIa0Ag+0Rcb+ovJQX5mWGILVm1xwm7gwMcQ0MlN1PX5nnmYGriChdvDHOUj1qEF
7vH3hiyzv6/f3BkyODJXTruJyaoJ/XuYqt2M7Ks/2KKHzXAGgshnmWy0DHICtQrYrc55xUW+VAvj
ESYNHfqfv2wH6iRDVoXPloiP+FmtSQFovSSqNiO/Tk2X/IBY1QrItTWUw9zQ4hvXiAfP6ttKJsb8
JuxzsdZ0v4wmyLVr57kbxWLuig6erLRx0Nvh+1LMXlr0sMmhcK29K+ISKZffhoOoetGJ+gpjAkl/
9QDdnndD6V+HmP9xJIjoUDb8RfEjuVxaINFJuAaDFUcRQMMTiEeCU5jP3IV1KKIpt92z4xNLYrFM
hGU7sEI++HDFgXwm6Q8Za/0LsXLnMeq1Te/I7gVMlp8OIYzyVsw4xHwTsbbiWnnSJOvbrhRyDrrv
oObqeyB7bgJ/8y5KRNjhECAbiiji9Ak42yVOArHfJnsb8tXhgZ7N6wpBU0QntvhfrDnwtsy/OE4k
MrWXjpWKbBX+5KCjw+o8PXke96l2WJGMrRYwtj3UIfp30JUtBdsqB4BMwtDh8kYm6NhwLByJDOUZ
k6d31Cu53h0iQSp2oX+CliO/wBZb6yNf7u7j83Nmi3efCUfdmjZQg6dLAB7MyodSdx5M19zVUiga
+cDLDr+yTzIvnx301fK5Ysifosuwb8KsDQekXdC7xOf6q282sa2oOLv8HA+mBgq2Grr56hLrauof
lZU6oyyEKjVTC0j0fwN8Z28UO2LckVdAmoQpoZTj9UJqsyo2C1l1q3NFtcIYyLnVSzJELammGw2y
Gsh5mtXrBCxaulEdR/8s1h3/zGM0+Uf+0Epl9tlBOrIACBklUF9DHebyrwQ8ImuhzyxLCRaCBUgh
Xf1VoRPz3EcFX3HLLqt1GOfFL1OVrjLDEUTTbVg+avtHphbKgsZqpxoeHjjafU7JwtQsW1ekXeug
5Bou49bMYhgiZa1mWdlr3rxdSIa0bKDPGKnPiNQBNhs74EwDnpnZJpcJv4J9WkQZVcD1uprMb5Ix
LryHS388FraTWBYvejUuHlJu2pKeaWbWlrJ6TxrPrdJoFuURT+23sEIpMInvBoyjD26VDnBuIbSE
pjW1R55nGK0xIeLHojdwvwRp6jPPl1he8jN95KM839n7Tl9KLKxl4NCP4gl1XaJMFRc0KfjXmNJk
cJcQTOYCIunrTZbjaJL3Hs1m1N83jnfO5etQIbtYBaw/OM9OL13eGJg5ry7IWALyFNyyyVsIZBdO
DRUweHlRNZ6Fdh83pfDJMW9kUDufienpw1VWOmt74PVCpIrs2ykCRmWPaa8r+b6/qcaB9+w+2gSE
aWGT6jAjEV3aK01IliKaIj2Yj51onCF2z0ObWJ6P6CYlrKuhR2fuhkumih5zNcdHfpwdw+VyoQh8
BG7zUjgxxi9gTN+DYGwwm9qESxlUKoVmGAUAfo01+h07kLshI2T2IRVZZc6NiKyMqo6AXTK8LaYQ
PVs81cS3fL37m7/W29qF7u4nXHC9ZTqYYXERC+zX14A5cQc0jp2n6gPKnNuBrgaI2yccLcJzf22/
NG/RNlrqDgW99kSL5XnbJZZMhdc3wUIi2YEj0OswBSkpUWWIwCD54zPH/Gs1f9iTipQ7ILf7imkn
quIHpWZtG59FPyO/ZiG7HFqIOoPEXbvi6ykK23przpVxrZsouuAEG7BDrpGRgMuVe4puQC6f+KIu
xsGkcvBeIddu8fzX7fyBasXp2DTZUc67XU/cHgYM3Udrwo3PL/7/0W/H2Fvj1jenerOR5efVxZXh
vWJiDYKCklpK8PFXNy+PePnGz9M4ZiFa6KKIR43YuhGp/DjMYh7o3gvD5l3vY0EPFumPV+7Bd9RL
orYCCFcTKm4KjPdlioLic3G90XtLXwqYxu0+RPvGapKFaEO0LzGquzm6XQATSjy+WYLh9L+0RwOc
N9/M9H979usy+IzfRRlsGg56nu/3Y+ovb7UvS+IKOLKccIWH3QoG012nxpaDVJhUur7tFUBhynjU
Wa9Pi7y7tAe7LtisppYZV4yFIMkEtW9ZOhyTZ9pp63+uOePYkmp0AG0u12pS5OwhbsZB/mnXyFjc
PdpDkY4a+4Jir6esJ8naE6HJPY0Yn5KB2NrpMA3lMAFOxQAb8Z1lgsW5IW8U4y6EoLj1/I5KFH3t
OiFY0ivfQzvr5lpUma8j8xhR+Sjza7czgI2c5sfZC5DSZ3PgAjKmk4KVSLk4d27ELgQDLikvu1vr
urZ7oHiTXCtZY/wdENEvcrMXyCaK6NtzW+yiJwtcKCqoDu2vJWh5NYPM6oJzGj1RCZ7DGfJYRszb
kP4x82PH4hwDZy1+PhBTR3d4mzN+fTmzIm1mTIrgD0HJQTQFJhys0gfsqajfvG5QAFuYoNjle0rD
wlup9Fz8s2b98xdsIQbsUil9vmHS7aQCK46kda9IEb6yOLbuSg/E5P2xbZ7ldU4KGHlea0gkMrq+
aZXTL1RjBkd9ZSmbXQjXYUEl3UUt5rG0B3BNZPvKenzKeC0q7w+w27MkEXGW2hVebeNGHTDS7jZ/
mcpu1ErdZY5hQ4dcriDgaciFODePXvG/UyaE5JZNvb389q4z9+P5d7BV0wGHyBgGATvRMImV0RGa
U0TnaLqwMGaf9bXKbnS4dZup/ejTQ9oSkf0suBjvKfrfvv7Ugnp0ilTDeKi2SmJLmOYD4VXUC0ig
Oiu8EhzyQxInic1nucYrgv/EgDcGOVnstGvhzacIVIqUnDQgm/8vSlJWDkWfdwUKhdoDzU3CwwR2
jxohdXpIcRAxzV4Oji9AE/329iLGEH7vxihMxcFex7u3FaCpcK16oiR+L5gtyNHrtd6IvTWeNY+F
SIEZ0BUqmc/hY0qrgXTX9GlQSDPCiBRbcP5NytE6NggW3LC9D6Bb2x8JqaGs0NQK2CYTz5ZNvQuL
LGeWPORpP3spSfCDD1GBWoc3Fp7vmIxwZsCDo4VdyCer1ARYvNmrDga93X9uw73wK9Y+wMcFSH+j
oIdHopHmXnONlpdFCPOr8Ldg3jTFWsgEe2YAlp9U0QqA64YdmstonYkJEoSUg5vhtbqq6eoozFw2
B3MBbzZHpKfSK51OjBEKZ+PQ4xI0YL/DhWxzHlVUI02kujATuq7heRStJvQxVIcoIYUx1BLiXDZ2
LSziADXB9YnovYRtNmOFZhXJY2sWp0v3xVUMkX/EyqEeCC//Hi0ey5iKM6S7Q69DDD1N+kDGvrOz
DdjAdRTkvE6RvV3FU5KRiZeGSkQZz5Wl7WOHbH32EsPxPlPqqeI02rmI9/2KF60AAov4uYQs44e2
q2wETbjG5TlDdYEtGpbYqx6ygNIBImImOTLAMEZ8eY7I7AGRPwoLRXUPKsWXCCuxwaL5zwFm/H2K
U92jxob+zq3PYGdCuYMBKgfkT47fZxrtMav6Ddfa2oMXcEA7UqfUelD9sB9i+ZoZgyXRuuQgIWPO
qq3tJSVlgZXO5ordD7fc7d4HUBZY0tZVqcND3CktNrB7WjAR3VaBuM6UZ83703Vt9DYA6ad4pCPU
RwyxaVCkjDE+wl1qW8yzH8XEKlTgj/luQac3CNMqCfgC6Zb9t2UH/x+OBOQM9nIzF+G8gEnStsVl
aLZKWCHjqhy+/FwV/MaSZrmsf5jjOjT5qtf+CKSf64KGufgcq3KOY61Rb0hBvbborD1x7LNN0zfC
+RK3paBInZxLUvXYRCuClGaxFuoxLsvw4PK4RUbLEd1t4LPB/JYl97VGt8sWD9scuyTWafpGgkRX
YgtQgXTd44l8b1m6ZahuzFykWuO7OiGoPr1PoRuSVeCQf7U1APx/2nbDleGO33rP2+tBuNFiqBBo
FOy5yOZHvSrCIoJZm4cCLOqYJyvPkohO5wg8qUG/qiCB+Qi8tQI+yTt7VkUkwkPrwxT7llJyK7zv
OOi9QELwwHB9MCMgjEAwcnmO2TXWR7ORAUZ3mmUOmJpwYUU1z+1GiQhbCjoX8/Yt8TQE0phDrrDw
Zjn8fz9bG7hetfX73/3WERG4b2S2r4hsdmOdzA/pyalZV7i7O0OilajIKZ/jcRJaOGh28q0jdel5
LD8G55g1UYD8qXOanpj2GBX56DsDlDVdDfd69cUP8UXAyHRP/2RNmWQftZ6hzzUwiZ7Y0JZD48Vs
j5fUKNPvFubXhkSkzpWP85+u9Q6pD1JOVTQNthXX7ReH51zN1LlEULw1u0h4i6yloZhCS/qBspxn
nVoZGdckLtdmHDBV/34j/km4E3uLDE/bfnzGEhcMXwK7Hl0TKbmyTRwNXQRjIXXMAHWM+EQ9M350
YU33tv16NlxGTDl1vh58oHDfWJYrhhY/fJ4RtP9w+kS7j827RqwoQf4HnOfqbjg/in9RQRAF3FVw
6V7LxiK5R9Yt9l0jn44wLzspOsEIXvxxoda46r9gnQeUCDkuEeITfAEOW8lkGrFQNmy8v9dzOMwi
jfl1h/bwOu0NxnZdDNrheNq2rpCzzGG1lSp3ZQ5/8efIdDESEUYNMVDzEzVAFTQ4TJRENYsmwGD7
RIFe4Pf6Y9s7txGcrXQ0Y1fNWDy7Uk6/SGh45e8kIoammIMjJPSp7eWe3/HuWPC/yx2/qmYOeqE4
ElS+k9SIan/4WL5yRhHzQmx8jQjQGAJnxgFnj+QlH6TX7VZgeorb9sadv8C0VmeNu8Vud04TKhpo
qb+t8b1sdM3TDrbXFtLNYQgrjJkr0/SdzHKVe3H2imfjQh/7waZYLEvfJdw2YNoHkUQAPOnxHTGJ
225Pgf6HBb65j33RihnYxwXFT3JojG+Wp2D4OF2omW4bbrvW+OV80u/VSJbm++T83Vidf4CAX8go
QFe5JDPzBVMgOW/cdRzzCOUPU5elc9BjOyF/zdSt3ho4ZympjuKxyalRZxsKVH2VgDads9VVwDvC
USIkL+CmqagxvruJhJvdhXuj2UzpDFI9Dz3+p78b3omPPIPvqT+LobI+qnhijyFBjRC0pGMn4uqm
ipG+6a0j+oTtDG9EDRvvQXwHNjN+E56BePdlBQ0EZPQkJFkY8FD5orSi8uojatxYJBJ63qJ7lss1
RQT1dSzW5lodE2aSITrfzM2B1k9n4icSrAIUNSYjwg3Ze1NJeduei9sQusZ1GbcJqy/Eyz6DU6+Q
0jEF+4FYtT5O9Ix8DVmvA//z5vVeeTrjrHn4FRnf/ufcUaXPFxLlFsSil8CGWupvCsupMnqAe35/
KWoQTu83Z/70Ws8haNxcV5L+uoejLrhs1XvilVvcEwmWpOqDFyKgC2hnM1uWO3K6xMtOsr7fNdMC
KygqeIo6y8OZgSFMltnQsGxAq1v34xd+yffcfIhWsjUoxGNtYA/EuEgI11NBh7I8Vq68kzpqFi7o
rMSQOodD9taFwIdSBGdeSLjjUJpNMWmS+Bux4d18de0iJzb0KICSmQ4XwH7ljpSS62scEGoh/Eyg
4DxbQ1AKlDl2rcGI+3aPWo4X9x6kvN8XoOhnJB+Xk2C4oYyY0MrUZt5U4d8sp2QxmDkz3+gRomlJ
eIvjugpOSYo6vT03YKb8CIBS3SZSMpR5vUCLhMzooCQsEFQMV6bwzEOMAaGoUVy67v/aZHqvqzsJ
04V3zkuWk9QKrN2Nzck6RrC+DCVcp+dUVuVMwsNGAru2qUiPNhb2C47VS1DzHHOYaeLGUvKBEZP+
GF/Q0BRj/tgqaakfU6e00EVcnC/hWHHy9924MmOrgpfnzTOM3GUI7nMfXjR62qf6xoTq83LE7VdB
I0bxUc79AsAmnHVeOFxXWgJomgqAPrQplEsdHr14odI+VOvZiQBfJNxY9N290g9qykjiLblQ8GEo
+j5oYfR9G3wfh8GWQ5fCxKlZ1gGIH5VvmxOm/ZKgTACJC89xwPCLMy4VmLBxZcTHp5xAhj2VNatg
j99lULYZqF8v9iGzsUz7g1VWPMlOfMmPhHHBRbGn5nbzXJw3I74bnK+SOmtuSxTCbC/P8vqIQZIW
5e07x2hp4mmbhE/6XEsIHgOB8Rc36hiJo6hWYULNo/fc6BYVcwoQr06ywNSM0UHl/4+o/H2BNi92
oGkCClfWfSkVkveJbPnRGAk6WpjfZIhERURkew6eJGM+DBGPdxO/IpuSRM2HFd2avvhwQkjGGWZe
K8B0q7s3pmfoXpJuzmkj+W0qkMfKEHumJIoTKWGkW5qXYN6qEUsrP/a31AlRKZazJwmuNUvdiR2J
FlVxc3XQsVHLixNWvE7wO+iFovjFaNI5QxIbL9YZD1IG92E6srTpf03TOKwiLiI+ARZwcmYW4E0K
KC9ETDlLEI8PGq4PwLonzv1RuNnHj1pC1kPBL2h4QFmBQOVcxQ+6QV/SkWNaU+1iFrI/wvH058lu
7eDBkeYLdio1b4sjS93JNSpGEBh6FhEG72M08ISdVTOYnwHJvPG6CpiMToAYgeMSjE8TOw6Co1TI
ZmXpAczhFGI3yn6H0JTqXp0kwLtWrcUUnE8krMlNhh2zwtJxMdi9UP2eakYRhhAIF8diVN5i7gFp
lcUnDvgBC5R2A7grRdyUuIuRzHoZHd/r8gj1OB48Bmop6WqXLJymb8p9JYxq+bHJGDhdkkqiRAZ8
sfFTOaZW/TMA+JQyLXYQejmuxbHmmvaWw8AFqBwLO6OKXXaclIFU6YwbbMJ5AWDsK09gOJ1BFVlU
O2FC7H3VxFCNkG+30EkP523I+Q0hvb7EsSViY4nJhMobp7QraQ0Sz6SUpllNVeirDWdsqeC0qUqJ
0VQrhOlIG7Bm56xSh7gjx4y6xl8v5kYHhiNK63qS8rF7IgwEYiy/u9/eHJgTvmyJCOUKLy8y3yKr
XIA27pt8CXaEn1sYBV+VOw5wKpGRtNAdmwFqOm/Oipmi18+cI1VxYuzwkEiJDHgK6mJZ+SCG5+lC
k0pTXcRSoUm36YBniJfkPiaiZILWUwnKQ2Lw9aKjZhP6XSA38jEyTAglneUK2Nz5rXp0olkaP1QC
aCjafGfjujhHIpkuH6bz4hzqKVoOqS1x9rDnqYwLwtkbBvD+Y8/ny7mBYJKJ4TcWI/RQ8rY844IT
N1DScupTOw8he9LaR62TQhOUwrbgUuh5zKF3L2OhS5kuHAI01bppiZWJ9kFuMTfiq0toOc1RhNk4
EKNlhKqbKquCMfPuURWtmbt/RsIbfNP8afCrUHtsFSWbmY7/iSIFBA+kBk/zJATf5TZzp2pEpUzh
Y6N0sY8IhwaqpiXkVqaISUgnPq/nGvKN6qIHmX1aFn3htHyaSM3LtgLXII0u0jSMk19xNEf9FL8h
IKPgqtyMRblGlRYOzFKWLySWHf72x6v/x9BMcYWfqTn7dGw39aNxwsA/tR9hjejcFxEhGcbdsncI
hlutSXHtoXBsEAYvhvKG4puQVkd8qfH7XpkcLCb/GY5VEArsJadmVl9aIJAc+Uw/+QH/97zyfEsH
v9t6h4F8yh+I9565vO/zU9Ot/hSe8CX9+pUDzpg9gLQK6T55EGaW6cQnR6r+eZN7AxWi4VQvPRMB
ImZ6t9pEjVZKXdYYcILHstmm8RkbFZ2CgLxJsUOEYPn+EtHhIjAVytmecxyuPU01EmN0a0lNEZyN
TSsg8AV6u/FSHKah1lj/us7jeFcZVDxqyFjee9+LoIP9uQM1Uz0DrWEhm2sYuLs57pT72c7PsDyJ
hrIusjMN9ZqUC+DpWHbehQYTXgMuBgpvmopakoAGGjfWvDYLd2rlrpCt5csiFXPVhLycR/11AbTA
tA6mLBPD6W8NpQJyy26TXC3EbFZTpKHn7FGO+6JOPoypkIevwFV+Dsmw1/fRrgePxAomTL72QfJJ
yQu6xw3Az3jIMkkiOINcV4HT6zWyhL/s/Ooq2EafgJ1L3QOtH7t6FsnNsFU2ENt1b4pXtPUzSNVM
73vLJfrhvGKl4Bu+JAbZJFiVUoqpNmtfAluZcQiwsZZhlvkwL10lywmNYZAI3LdjhHMussP40Jiz
MHvJ1gkv8UXJgpC1bikA7XdFtxvLcgQmKTQACZ8SBmE3j5rIDYf34q9CsqXJt/IOSaisRyMwioWO
b5RCYh57ZT8AqD4xsk/uVvxFpv8uz01dhb97kcC2TncyVOxVF8qYZuKvRle8hy3aPerurCyeq5kF
EDYcANjHeaGeGvsevyQY7MpYNEXLAXCEuwmxoppwyeDtFSb+U7Nbl2nLVPHj4ktAh62hXR7QHOIj
Yxd8I/hetHZ6UPYTtb+tjvUyAfSfFxmw0BWp9UB+Qy+ztqRQ6MnS5f+kB92u/4GPMwOd84c9/Kb7
iEkQrGbSrdc3uVNpaSghCtDLSQqskjW2qOoz1pq9ZMTg5bFkgzyke0H3Ct8Q1IoLcwudbWvJ0pqw
BTsWteeVQlpPxC3UMFpvf3GfW9IXLmtofpSMTIvkdXQe08Til2tLC4zYEpMEfbM9eizjSd7E2ud9
+gHGPvFT9wzPU/+oIlO+awbjcbxv+CxlhFmyGrRWXEoYoKU9CnG1xUS8/+XSTX6ArG/hnHN4hR8j
WuD1/n71lxPO4I4KQdIm5u8extW2AKq26Ugvu0JvJbw8QJlUpa3ka+GjsbW7YIvSs0W+ojV0K2JD
ps2RzsOktIEMFp9r50k/br4vD6kwRX5S9paTn5zFK5041Mf0HxDviHmnyjmFvVzjKVVqsvyWZWol
en1SduehtzBglTJyFYPhe1r+njAiXm2S8Sj8UOmm+z3DuggRGh/6MZgh3JUBx2QGYJWNFvzSK4lL
a1wsagKRajuuvAiGsLDECwUGsaa3V07lsElAfPkOIWOsk1bLyoI5Tu6ZdLKTuV2XNPYVXyhLhOWp
AMgvE0+moxhV9EV8r17kFiyY5owlc+yEbEkeXgxvnj+6BigK/H+BT+i5ncDE0PA6fFIJmztblINa
Rapt2TwSGEKoQX/ROkbyhM9Vp3GO4HmuTthnXO0WNrO9oBW/Eaa9dBn98iCZTGQN7NdPu+SNs4mt
O4jya5SYZWvfbQfcciJXZiyOSCtHwEEaL5h/vQLUc1ADZuBkrGCjlYJXuhNO1ZK9aB257hUSAANq
ni5zeeR2+at5NMzFRzG+aipX9G1nlogiGYy/xcHLL7Hw7AWg23nrweR9OGCSrMTuVviMyItTTcm3
UuMvS8KM+9n5H5lky1VWfAJIQu2fFyj70prmJjIG7b4yI9xDZUDtt/a+pxEKSomP95Lp/AePJzNw
HbTYuxPxoAF20tmQqTjiTYeEX7LsxUdVw7l74rwjVvVD45h5egyncLMKwY96vZpGQEO///F30lLX
8R/ddcuxSHJJIdXrB5Ormm5HXmtHbhV4SXWEUTKOiW2LbqfwoSYfGf59IytixTEl5TrEEPEt/ndJ
zcuYy8OgD8MKI2j73nDHpndxJpym31vvvOjBlRskRbDukyg70wIkr1Cx0rXtxdzLESPcttsLMyT1
ufAsDIRU5TYHhezndnncYg5oF4VvfRvsJHWrXPYBs1rAN1aTPngOV0leWH26ELHuZpZBYU+kjeOr
ywmvtgDgMpQa/k6st0Vo3TvENN/XEIl40IXZtZ0bSs2UvZ8H1T1+UBBB/yPbHMbYFKHeHEUxfWxm
/+INoIyiGnK/5ympuIN9FXI8NMn91BHe/lt/SJ/5Ux8ETZ3sJ9TzDMQoX2iZwzSbrPMMZUhrB9xe
pOwyLP1PuGc31obRpooUZZLoZIA0vhnohkBrZBcgtAYY1obg8veL/LaKVjQvdZbsWqBFL9bp5AOi
Avlon/u+Oz7DBfFLLWjiKsD1Ymv6C9a8EjKHMJMYeh8Jp+Rdkjj/wlOIGoadza+C+Ond/co5lzlK
0ZYvsNzZX5nlP0aNrbuqqaDEykITmOcv8FUoO1+cw/maK76qMjLMtmzuX5sZJkl1b5A8Evc09oQ+
PNiqGMgrWkSEazjg7/0vg+IglVD6/4Olnx8gt7pvjONHTyzSEAwRaJPeN7LBoMh0DxBt4Kpqw/mz
OGLyJEvQJfQJ8QsaDS0nRbH32SWgmkMYlgWgQF+lmwzBrTaA7hmGQKdiEVk1i7hskhhlQhbPymFW
FjQZiQLXHUG4u+5rh1HVdGPXBva3Dkflpc25WqRAtZp9fKI5+gIdVc86kXQwf4If9FO1P6bYgJGe
kSGlDMaCzP8V+/7NDKY+iWR9ZTu1gy0Bz7TtgNwYHZ1TE8hH8zSjCypHRLCST9hCgGux3JUQOTVg
v/RgTc69wptJNGg9n6jzySyhsOVZzOuisTVg9Ami6FTq4qeEO2FI3hytlRZQOjkUShmxvldzvTGh
cBBxXhqo5WHA5dGVrpMBi5bZOwVWCStN73ESKgHBnZObZ51VZWKxgcJB8jrID/fBTNW7fW8Te2Jh
osExQullUvbnKtxur2WGTcABYZyYqGR/jeY1xyUiomiSNFHpnnf6iICrFI5B4bHxZq+OHgIP7kWy
i7jDzxJ5RVFQ4pRZHQ+0vULIrfEGJ2AJrcVp5yL0HPBvJGu4piB8+9GdvMN7SLmT4fZ4iZ2h4KtM
wedClOc5c5QXaUgwCVs8Oy0BYx3doYeOyEDLSelKRYCnMBXSRtnUAs0JjdZp4OXcmgRe4Dym9yeC
RTCTBJGfa3nreFUAzQ4v1p1gXCCfm84OpzMfDQeSqoC/b2VEm/IcbghOKP0fNOsWWk5XAht4CeZh
fifi5ZlOGy9UrPUxFcYlMKq6g5rKbX3N+27Cx5q4PJjeBqvayT7scCPTBPCEGQ4VjmNoj+SdjpMu
nqagOclec78ToOZpEPkG5PsSf30kbUc2E5oO/2BCz3XOyv14fxtfrjLIBkb8JoFqIL59lMWwgcxF
0BFxbIYpbDbMiL6wV/PTu5xyROUzD5MfDVellKuY2Epnxl7NG2rGEY2JBlPWoL7woPHKNI9rFRhE
Q8mchb7/qtkMw+FSle1wiSr1zDSx1bsqGc9DbXhj4vXsEuKf5Qsuml/3jiMdcGLUgMHiEVw0EqFP
LMbTGnrlfdbN4WcvPlz7SL+FwxmQQxymbQegPyQYzdqLWDqLBrgLV2MSvMJIi42mtQgoN3dIxIpZ
/sqN9WW3kinYMX9hzp54KW1o34jsc7mwP0w/54O3m9GdsnnEhjKYLER9Lg6fXoW7ZOyyEOcuRMJe
+7y/zWe/5FP6NJAeqLjsRq7DbrspGBn5zmsaYAFrfThAaVWlyfL8Wkh+1Pfb/OBP11QECAK0vRgR
/o0Z3alNl/0tAmbbuhJerpKIgiw/WlS9hMNAltvh4ozGDO+KJNxMA59HwXKwah2HAELZ0cGLejbi
YpxUyCLPYHwrGfC1bokNO7FXcMc7mvMXqGagtI3U1jnppF13X21tK7FKKxCqh3+CmYO6rjbiwP1f
dqdAghfB7SBxgr1vh0MXqh3km/dEqUjNJcvY2NVxA8U6x8/m7hzKs1cLZl0gV1JT3A6vho3gnWkU
Zsvaz3p02ctJau1eWhEhbTeGoUoEN1SkAmANsDIkuPbeLEhP+Ihlqb+JNHb4L1eN+z8dvkO7QvdS
XFbDW2uBMih1dVvmS3Yr4My9aALYOI+uHUAHWoeqzJ2LYzM0HAHjSZWdyLYBGX5eK6hpU4WVbzfn
abmMln2FAdvJt5RwrNaLMeG3PNNCEpPak52hYqxwpuY66Fihe9P1ZhTjzyn5BDdBC0AdfhCMK7P+
Xv8PzWIUlYWoLNXugQ9yWwHOFV0LxqyLMHg6HOtptO0VxiLXpmyprRzU4BJNybUzz4j5ehuvchGB
/AaCCo8Y5F9S/9eFu7jVkeOJ3KI863wX9X636P3VsOpliDuCzhkZENYFQ2yvttrp1Ydo1l3HgOeg
ZlTWsmR0OfwoUPqvZYJ9MT+VQcYSMUfPNYZYHXyT0w4ihUgx5AY0W9kLCTXgSaYPkpvOVM/KyzhT
PRQuLQwhNpSCCTmyEa+KwphaEC3IUwKV58dqw9FXfDcfWk0S3Q4OBstmLqNyUg7bZnaj1SaSkhDV
2eANDRzHWo83m3VIPcMrPsxOoqTUMigDtkQ4UV4ekIfMJZk+G9/M4lGY9dfhYc+DH4uJhsMH1nBz
AA86IF7i7w7SF+w3HiC7KM/PY1espzdiHFlUE3uRcOj41wBlyW0VOqzBH9jmN1DUtOIdyG1yn/94
FN6qnZO/7ZlM0D3Sjpr2s43i4vVhZfdZOLdvCxy8EtKY7zU11vfGLuRZ+bP3rCk/4cKKPwY/eu5y
wb4hxQVjEKpHhKK1RH0UZ9TzETp0OOMkoQO4mW3rrmzjmhb3qvz4nXt5LqM2i1Gb1Uore9fNjzsT
x+rq5cphLzaH1oCu5swnAdvPtg246IToAnzo58BBkmyUui2+hXT8oIG4UvRUS1GwxLgVdzw9TRBS
hUDQn62Qrq4R4XetEZy6mmcjCTH6UNCGp5hemwYHeS1mWHBMYIX0WT/sUIKI2f5LlNjlY2ya6FRp
ocrIgLQQiib3tKsGtD+F27yTVm1BGXPoboZgCNpenRs8m7nJbFsxLKgltsLj0FAQ/O7H8AQBYkhT
Dql44/dUCnoW1KsHudHRyDErPRH42fdp80w7UqETHeWmEYLq/rHQAaxJvwgHGb+q9aKtWF7eFZ/8
IrcJahn6T0XpjuI3jKzPg9PHxw6+8g2C04HFiZ8eB5Mk+owYis5tLMNiYQlmkLV5NTpzJ77dwu5Y
TYtueejEOigDMF/hjziVd9iIF0uVQgB3V6q9c5PyNJNcEQCs9Wc3d903RpZ4PugUWctENGbJ+6Ey
bDn/BBPvPQfjLob+smLldBjYqhmH2gfUY5Jw74MtwOq0cGlqj51377KCrK5CouGluAYF6E1Ad/Se
TqFmWZupw1Fld5nH83WnDvdI0lH1GlOM91MhPzRYF9YEFDRjDvmYXUakZDWd7TwjiXs9rhjPeFBi
DXu4XqAv6LxclSqigzZSQ92uLxUA/5Q4dmfCDfEq8ykGwbfYfpR6lwJKEOfCNzW/XEW6vJs1Xa8F
wfWDWqkCO7T81v5tEz67Jp9D3f5RcuYA3tXGvTj2UxoVsqbhuS4lhi8+swoATI4pxmqIU/Ft3jv0
CrTZnZQQPE2XhJD3bZhwSDUo8VG5Ar/Wm+SRxeERL+QqzTtuFwtFTCgZk2mlbUN7XD7mZcPC0+Mv
Knke28K9JXAbRrsYuQCzHGe/Lh1TwDM+ELI97EyaxwhBsvmsZ9QTUPdu+l44NbDTsctUPpbkuSar
73+o1v1Yp4My4PBZEyq0jmhR68z6wONL94SwgXuddCmcRDR5R337F4KYfT+omJeSF4vAmOgWXiGi
Q+71QN/Lt8kvVIttyVOpZCrRC6yHa9bmJfNWVv+le6rQTlO+8Jdic43GOgUloUGdt5KqEi1+L2Ng
lhhMfHYXmf9uEt+Vb1w0vxahe84FXrgCRPxebRMYONdJAcORuMriFPZE//NIEOzDpnzfs4lT6GXg
MdvB0jdLnsD3VqN2PwpiFzbEdw/LzNi3qYJEAh3SxwESdrM1ctEgPsSNnAOWiaMo/Mmzoj4s73MG
WajMsK5YCa9CBRop9lFefe4de8J/DidNzObxC+vPu6bV/lbV4XVG4ER3BHjEPsgXoFngnDPllQwJ
rQFU54B8J+l/k+eTwMPSNiHDm9Bw1HXDHKM5PSlpWvfyQadW90a7ndk60UmNAF5I7nyc9ajwbLRb
DdgiuencQLDTWudZUTVBv7IAhwXgREfuyqSzKwfcJMC7+OPrhn2wPDQMulYX1GC0Kk/3Mj9/8fQi
zrwGAMBv9iugkzAbzsa9Oldnt0dw7DoubPjA0lfprCjAUcLURwTwegPek8XuZ7dw2QAYTqvj219S
xVim62/0S+WRbDdCOHxUbXcLr7WUgeyY+ggQs0plOVO8SM7kYpsIDHzRyOYRZaecGAWdHqhdz+xK
q/3WvU6hg+nKdxhtuIYgZW5mLvOiEX8/y4iU/Oidb9zCxpV7AtJ5NmTJjqVrM90jDklSdnpjoSfE
oTkIbEZHcXORe0+iUXWCgqL9L4YNHcNBu/89cBAekq+vvaKg4IZxKkMJOLOmg6/e7jSbmDsOFYuX
Whu2tWQda+BxFLeySKUEJCnvkPgSupBgj+cSh3N8gy55CCZlkW0Tzdgtpe+u+38rxFO/1u3Hg7Et
V4kiTJMioswplHv6+O3T/6wS95+cu7yLkpT5w0Hc/cUV8Xxhud7vy65ZJBgNIHMVV9yjuzo5zAsF
Kd0YJ9jlIO3qM3KCPDE+r8ufBPHsb3TuY2lkLVtO/evv3RJ+0bPJi68vcP0mlFJ6Ah25tRExG548
EWkzDy31yaFZ08kYUGT0GDUVn/ii0YB9yPgPI7upHKPJL2H2CLZoDI6Q2yPswDmAb1O+HQrUVhCq
TJ0idpJNdTLT7kbnrfAFQWrMoYbiiyLOY+Wx5SY7VPtNbaCxGq6bGMh92Xq6LUDOElNkXsfhKSxR
fNVbb2QP7votcKiikrXZjbKtN4QxMgJlhggN/vFDdy+b0XLS19TWRMrwcsNyY2X0Lj+DBdpwkj1A
5r851XlxEcK6iYibUIAymrGCSFh3QivjuKgvA7XHR9PbGv0Wrr2/qWGZ5RlE+7J+g2LpZ061ZCul
G6fWzXJJxOoibdFq6a/UZigP70y0X+lqWAvImiS2CyTxsB7jE1WuDrVuvoGYMmtDlWgAbYNkcGKq
RHcE+3qrpRq+J+zjQ558JtwItYZYt+Q4tQek7OTQrcHlEthg0R/YlhWbcHghwRCIQkzCCEBmdqCf
xeM29SKmBEwDJEfemQMK7OD347MYfqyMdoRmX47ZbqJuTqQgpxIwd1Xtp9wSyZxDEQ194LLPkLv0
BxLPejVrU/YUfefKWqva4nbjcvk3juSMrh8SKL5BaBOGYpHzTKQKgYejdE56Kve9wpdU4nwvc2FK
Zf7kXRx2dvbxaPN3oeROSbMvzZKHJnTDcuTNbc14o3xLdqCrxBJ1qYu1RHMivLliLFShDcmRjnVE
FVn9g7RqkTat9Ca/tmL4CYn1E3VNqtOpohnOtG7uJWB2PlSNTq0COyaglhn3R3X5mqCDovfErEzr
E8CCeB8N5r6MtKcVFNQ3hnI66DV5sxKT2Dff6I6PxiVVx9yWcr0JXQ66LBs+XbQYmRxn/p9nG/o8
3nw6PTogbZ8wN9BT2qpZiGzLOjBu2225Qv0LNCawRs0e5CymJ5vWGUmgA30sIbl7q+qp0au8y01K
fFpb8k6qzywnCCXwNHfie9aK0/cSu7/sVgDkE/NrlldpE4NgC6hlmse0CBgS4Sk7GixKIoi+7Chi
zJ/o4XerAF5YEkKCc66iAAmGhqlUbb/r0PKAnDvC7GfhVXMvNPtvXUrmTH28/YrQ5gcsK2RNovAU
QRhqxVuxch9HL/EY99aPRAjzMhc9Rrt5AkUMWRgZcwd/ieKZe8O9+6H6yinhAfSAmF1qgtG1wl/l
5TdEnGYD3YJaJjo6ZiAtBtq+raUzXtzOSwcs7do25HehJlpqkUpBKYaQyALeY/Nm1wyl0By2JDAb
U0xBuM0/07qKOWiR0qnIEusz4ted0Dd1LKNIRNlVuBHsE6fHnKNAUkNvjCiCBbzI4SUomS8njOF6
jwnRlka6+cV7NgXdizYA/hcWZggif7eUKMX1mrU8fv1yvaaXg7ikY5aa12dkKchwIBv4u5+Vpcac
BQZAq5Mk31gZjqEcP54i0ap45nnlcKLeIHTbiR42OsFKXZUgK/7Tc8WSaS9GFSpDEamSpahS9lIx
GYjc/Y8gQ4l/jypHIhGhE0+CPueybo8MWaE/gD8HyVyfhcTWSXh5jbi06D9YsNp5w1XY2k4/JW2E
BjwK75g2NgUX6PKRCJWqFooF1rJve8cdAJw1nZMpiddp5BtzKlCrzRowQReYpoFYZJ4h2HiUaBVw
iGz+oEseLuhri6IqUFkV+sH7TE44Tl9lfIV4lLC95BPMNdw4jv2ygwkobuEpVsjXQ2mvnVrI3Orr
BLhLJwjyGITvMC6XzeDiduaceZuIzeYJF4z3xMwCrvxL/0k9fYdkumZ0xQOWvC26zjY+7MvYSgEY
86VsXlNfrhTHWXNPO6BvYT3mUjOD9CvBXpPn1eFvkosUUaixivJAOuhZJQbj0FlIUt6jgpubaikZ
9gADfzm8QwP5uVW57Wof2ucLL0TxFKKAkPfrvEp2gWrJ10bTtuKghSEr23ea8gqOxCOgIh3JS/6+
GnMN3vQGhY735WrElKQfUzE+RhC7WGeIBYmQ/OJrdqpA2Pw1QtT/zYU+9thHDs4d7FF1VwIwbx4d
bU/lsb1G0mDHHJg/o8EmaR7Qu4FUvruKTIUcCEUdV9sgTXdqbJ/dkblRwQOuCbPz8dvwQWOZG/rm
v8/fF6QEZxV77yFWd5j4bjmPLj6Ngw/4tATnoYFPs7A6syOj93fsyLoK9nNxbldtDY8y0Su2pgpG
oyJL37U+SjWAV0LPmxQy+owA02ehB8ue1pkRAyPipF2wHQYbc7vf9SOlvrup9KCiP56TRPaNsRnp
Cz7+y8PcQMTBZRKL0ekou6EHD0e6X+1g8Z+JelOnlRYXL8/qYW8MRamBobIVaNXJ4D3UErpi4Blq
IjHntpr3/vYXXOXhuHxgyTGuNqR92p4X+YyL5U9FWGQAHqQU7EQb/39TOr9CErorwcOLZ4bMlk+c
803AUQeGvkKcYKkJV5MbaCYBW3jNSp2dfQDHWzzk5zYjq/fiTeCJOxBigUm6r/zpfAG21AUvZ4gk
DQsIKGk+YVTy0N+wd/CWYtTIjo0xKAndlHbylLGxjpTuEZA3OQrm6IC29n961/uxwJFsX77Ohxzi
cdKRw15KW8XAsNSrlB53GiTuSvuBBjODg6HsWUyLWjeblQT7pkXJj4TKyTJ84RPDpIDKN9KaQITO
0t8jq4b2R14/x/0DPlt6VkV7OFNCSOCNmRod5h0hV4Yfe+rMlDdxo7nQiBTppmXqmPaHU9lRJKzp
sZA8iUlZ2w1uPKYd4qEAE+tLfGpc5fCFfX/QofiuwdpZ4OHsDsdATkwDyloiwzhq/ZSkz6QkkdQA
WRYg+lTl1GkrHWxUlOLBXRvvCqxtk4pnnQwZ9rCsg7ezTcZxuFho8GSieXhgSeq8WvX3szHqhCQQ
B4Yi22EwAo5troIvmQq4/66gcINxMdgMY2DJqq2m8kW8J59u+59mNexA4N6yZTIxI0IpkR0G22bl
DGO2/JAvu2TLIdGoeaiWAQ7sTiM2lypphEf7x6P6jbw5q82U93o2QdBmn+Z5ZVZdDlkRxKoFl5uT
x8OGPsIkpOVdqHtbv3juSftY7ZqnwObC6O6ttdzjYu0oY0+tsFv/SaW7N1MReBDXMTzy8s06wKz9
gviMnIWyQtZlw875W4XFmMHZbmA9aRU/q7Fp+aeedExyOO8TnNb3+LADUvcB9Lkop4xFhlPfo2rn
V3EcvacwXDbH1NYBeX29+0FnkXAMRyCU12lKglGqIyXRKdijjMaWYKD6nzYKQvDoU58b8CGXsNoX
HVCCWqxW2vN4PTMrFf64pFfUhhOW6MRnoJf94OrRw+QwKPTLZ7Jh8G4tHuWE8NTgev39Ni3TRZzI
D1AAy4+7U0whenj2hxvWM0CD9oWEDRwYv/VW6ourIJbTpOkngXeqINTlwSrjukgD85Uk/pZGzlc8
msSZBW+Qah109R7QSFFhWObj6wQ27mMceZAjmEhNvkzeD8s8W7UM4aelL7UDcfay5d3CSNy0VxSr
QNGunsLjfpJOtIjwPexYTrv0uOgV2OT5RlKRh6NvPdeQTkxUnGPPKuRHaUoeqSlB1Ak+Xs7Iedn0
FxoG8mfwd+dVq06NHZEnsMxYER27cbspp8Qmeu+++BP2kBxRJC11jWPyoeU7ze4OVYfNOVVtQ8KD
S22wRnu7RHOEBzF4ApdsruMQmrXevbaTfqeo+EdXno8am0sW4McXwz7c4/7m+Xge13WgeJKO81/h
hN1RXqI2nyjWbCkP+WiV5BdlOezwSUjObIEed2MBwvMkAAdA1VRQcfcIE/gNNfzL5BmDLYr303QZ
LU7xCcZFlWBg0V325ubF2oFGRJpMILzb4U3YIeiHtjeOFwosFu9Ebk/wGYUNTJE4fT9aq6rQPP9K
B5laXbJZv7Hw6Y4ziUXH1HET9/FHf9XPcCyZuKw8azCqOXCvpSfPRDrHeZUnURo/zHWO6kcr28tI
mVLJOjjyBzL7Oq7vW3+Ysf8q5HmzS0EeBHnryk8CH3jKytt2t0Cam8fIF1KOpRLEvZbb55aQTlVe
vN86dvoPYApgiMI3z0Y4S1G110GYuRauDM7EfXrjLaWKza/ePIvuTb0JDVW4KZk4+4j27T9/cBme
+zSXeik2NIXKgoC/IsEiZ+6J4yBa7PAJ2Xuiulr9mM5WoiuA2onsd11iK7FY+XVTp170Xz8BfPDo
Vjm33vCP7rIYTCJdLteAVwvJ6nhovC+9hqdI4HH7tBWx4fpixMpLFMjBhsA/mJ2uiTUSrJgJGQvO
NqVNU8fCn27BtZshJBi1JdbnqTWKd5F4P/UPw3pGn5v6S+9OIsUY40LyUJFKc+HMwJlALfsJHfF5
TmANBrat7NiUf4JTp4vzLeBVHjrELLhBIsRNzEo45VsrHaRtmhASFfsH5yrK6kemTDCgGGTDR3nS
DmPGFOxf8xhBmqp4zs5krCCXyagZYMWeAvzVjy5OUW7VNBRHl+AoRL0fVw+aHPJ2fUCIMy1eWRZY
4gjO4gkM926lm0s81y13l6ssfziok+1u8l0oNARtmB/oV6A18MsW2geT8Vwt0YuypEXgMM/my0gT
eP6WtQd6/AJhWbViYlMH9+SmuZvv1ozB80rj1YssbGwVZ7QATqZwPC0faM/u0+3Gwg226fQA0Gwj
harwGQ5QH1f28zCd5jv6SKe8jSkJtA7G8gpvK4/tkPoWU1apjZvAhxuZk7ZezoxWSMMiL8efx3/h
jvT1OTxuxm4wMjBKHe3ntVLA3RSpIKzSB+VxOxEpO5zK+8VaFStH+DwthlDuBUPnBD9iB4esHfDn
RkxXMbIr8uNNTHXnlf/1mqaT5uevgcyZ+1ORgmOSA9K4Mkv6ZQepcnW0/n+XKknM5g1/fbKNfA0v
miVXHLuaWFOK9y86WKS0BSLTliiw2td4lVSGb7oNfGv+RO5jZq0uIKy72anX2pTAuAhos5Bm1Mi0
ljp0xsXqwYiTbbdIyiP+LPzVeOfUNJXtzihAc+oaIhi3ggXzpnEtYdRQp1SeBtMjPyX6sz1WLT1k
JSjajGspKghU9620AF8JQmGpIW1HH4EnV5L+uWaTStm88wQyYTg59f/0pOlsFU8UzErM+cZehwry
sbuI0JUKpXqc8C3gxSC706HpiwkVU2D9nvt/xkhdaAYGblkYXUfeseVOkXTj46Q7qkbdMEsNr/Oe
AcpDh7rWv+j/2ePpvA0RPB0d9UOVRnxfg6ByBdYikmb7TCva9Rddz+4iYT/265hArGidey4naZnk
eMqBKXhyzTzu6gbJ5HofgcQ+kIPsY9O1+auZD/dR2y+V9RM3WTNRTLG9I6vsO91VViU0k4N5CPjQ
CGVowE9kMbOiJeGlNaolM9EOQIz21fbgnJwalhrXenzEp4pxo6NAIrpljnlp57VEPtd7v0yxOJqK
mJvTw4I9Mo3xm0tkVMLSONxVrp++NbnsGWMKzNduYQsgqwmg0Ytfju/2Aw7qKmuvrwzhwFFpaoqV
2MEZ9K7Sx1lDJB3jv5yR/1WpCjMxDYCrk9zo012IElDna1nNxIubmgfWl9wOUH7kXPxnFRywri+F
znxlfHcPP229F7mpUqGDdvUk8TYatYIdaGZX4rATf2gHvIekzRx1trkLT5+gvIWJSeHC7cy+gtTX
gjP/DMqDf+/WcuD+y7WaPHYW0mprZAp73gNMH4fHlQx7b7madHaWrymRAnQK9HXxKwkCZBKggvZl
+c2eiEo8rxiI7qPy+SqYIoG5VOelsWyVAz+ppHTDM8qXtDAc8lnUUWPXcgy1IoAdU7H2+hrmpBi1
6rDXSILBxNTeQckA2lQNXrFcYC7hQ4IC5pIxbXB3uU0BlO9X6hDTqHRvoC0wCUKRNzrK6YaRF4vg
Ii1zFXNZFmjaYuhiArB2x8xZBM1SPI3qxWLqbvv67VbkFEhkNJhKHUJfbK90O5if7nORzPowoyPD
D3KCuEhbD+IY/nF5jkwb1ClKi6Mo4Yf+zBrxP4nlY+Pf4JZyuGA2umy3QvnFbzTwhjePeSW+TX16
Ki6VuG7yG3+YuKixABka1M99Em4Mo4L1BuAfPIkPL1Cx2fBxqkVBhYCQ5MDplHJJtgfEaKg4flDn
/WiSgoVARjKJvsP6RsnXoUVGv4WnHmz34ITtC2icgmDV2HGceJZSfN5oNttGg3EooDmOwa6IHGTW
CvZy7znfE6OWvBh8PYKOcrd4bJYnOqL8tAbMvgRNo0FYwfn43qIEcV48RXRO6jJ0DqmPkKlSvz4o
PsyWdCP/CwkJioKabJvg9xAANXxTtLGYCBFCgH18KeWWm3un1/u3Z6JZ1tH8tlP3WJU7w/HoC8O2
v8qG/HstaNYGGhAyKrh0DTAOjCgSM4riJNwRQZvroqfuG8t40JeLV/CYBG3NeF8tzau+lHidfFFB
IysK+lGZPDx75nPmExSfz9/Sn6KsbJeXMTH0FcX1kFcCy/1NCdp0Fzm3H81aEv1NqfcTKJs8y+wR
sDy+pNMnRavdBqaSdTzXw1nfpd1PoY72BprLiYMahK5P1KKUCcuouHyrWw1f7eBwSgI+KphfTFCh
ZCKdkdZDugxlXNohUaafaZRyMHnsm0pB90h1ge49yu8kmcSw0e3Fk3G3wKs5rUVySlkNJwZ1TWBK
4TAo+oMkWQr8KKxN+Z6HiU+nVlz2NTErMMT9fgCNZZBZ2R1Cbl873yIAc0MXaNkAeLr4vV4kKc8S
fuqZBBM6kC3ewn1zloAL6eqZmmexxMpWEdjV2gJ8vimirQD93XJ1zrgB4KCU45F+sGwrNLGNIMhd
XNtPEvEjL5UEEF+ArE+p89lGuAvTdhDPYBTT7755XPa7vYBOs7Wk70A+bmVoUt0Z4RU1Y52CGvhP
pw8PiyV0yxe6qAHAVtLMrNveLnQ8hpP6yFtMm6YhlF8Y9MM3UK9myUfuUqqjQwR+P50wqqgI9vg7
DVLNwoucXF7dZ82Px6CQ+4SH+t7XXz6MzI27J97KE0RfeMN4Gb9on4Wx2X3SsBN5cjxthNBxmqmb
za7cJOW0wsXwf0X6K7ww1BVdn0Isig6soPt9hT7Opbc/rZEbcuLUuCDSjCH0c7Pb7EMyaHFR9qqh
K9e5hVize+AvAANeZQd7ntmQD2QptDGmpIHeVbS73GrDhrCJxqmLy17Y+GIU1TsUjg5h8YdzX2Xc
yCC51+Kf9mDE4now+usWktPSbKlzowjsDNTWklKFEXZIu6s5CDxVAceVPpDB2q2wcVsDn+yqWy21
W3g3QV0W+MS9OC2vZnVCcd4rRSu9QEH41UA+BLwX0rVktiCnDI3XeDo0TLmFIkIYK6OWErBxCl3e
mD1Qo6Dkt9iG4pkPE1zubV1o73KX1ZjCtV2WJKywt0fAaZdvx20blwd+oAsBe2omzsqA1mfhpFJq
UtX6lN3JeooEWaLHnIAAfezmxeUsl1g/ufhpGH13evIotEJVYChd7DcD/A9iMpGfb1sE9rG36qqZ
HYjwrpbbQ8O/1B0OR2QzZe3/iJV1eBDxNRZ+x9z7xs5wdPEsnTMLgm5cgY17qUPMBFAAdor9mg/P
ZRHnSllVtG0z3o73zCGO7vyAlEAGroKpmXSybG8Onxx/PxYjkxe6sSVU/z9JB2cviKJSV16sqQ/E
1kquTr1WGqQS8P4xV/Up8Kqf6R6HotO4lsbEmO+Ne32P41/bcjRRF1Kmha2GWwNRoyqGVWivFNyG
OwOK3xom7smFQTUo6xJ/eTgYgYOFboIPj0Rr08Q+Tsdfe8+gqsX3F9iRJpoK6FpboyPYJGM51YiO
5f+3eGbfaQkEuD9ezztmEe/dCbRfHS5OBYErh4X1NTxk9xp+uv6lx4Yv8jHAA2PS1LFRqUoEO+pk
QV01nqayX310OFKzCU5gVILklf4oiZeUs9bNwroQq0nUhA+h62uIpOalb/3vI8ycTFQy5+rZnu4D
Z0+K13DFjj7kG3hCPvZqqASHao2DTG63lYueyzZ9a8G6RzLE7yS6jGbMq2BcEDcuLUnoRST8Arna
fJlKepYREZEDraCIKwpdFjnRT8mtin2gt/EODsDOB8BUWnDWZaRBfWHY/yVTQ03XX+ikgGFb2Abx
YxBEPeN80Me9MDaDItvrGuhRLfC9SItMgk8JqOn8evJM7lhBV7HQOVEaNr4KMXIWk6r5qA+eAtMO
fJkHtpLLjoBBF24kw6V3l/b+Dy/RcK6c0SCHfWFmNvgRAn1YsElXm0LFT9Uw5aX4bYfM4n6Uj9wp
U5HZe0w/hRbmPb4DXOAx36fY0N8Ia99UI3BKEnSl9hrwZnnhLnzUa4pjfl8hifVN7lirFR5wQjf/
A/MV/w+AZgaCTdJqRiTP6oGkx6at8LSfENVVPTyboN2SwzV6HBOAGDVqcpqbiE4KG9nbvgc5KuTx
zUviLcOIASAUi88VJUKLtsbfV/5QTv80GPWrmNPea2RGUeqz8FeKHXZzT1t7yWX0FSJsxutYv9ZS
5yBM4ZsDV7azCS/8+s0KXZD0+oI1ooujX5XfrLqSTupo7WE2TE8sAdU9CWHqMcAEf3Q/FcxAYFLR
lF0tZFibk7d+0emLzoNW2drRGkhZaYrIyZv7ZUDYpnnD+C30oOTD7dUDwfkwBwttW//BB0n22XXS
3TWrASpkDRsnzsjHRW4avsm5ZW357Jhy1FKG94t/qzLa9F99sUGtmskov14WbjqFoIKenGVXXzNV
KldLLD/5N30f92h+MrtR6U0YWZhuIWedIYKdn53T1I/JFttVwZQRmPk4gNLnG179O7BTUMlmQaXo
nqc/yXTLHvH/XOtSE+WfTb7zeVM+LgGhsV7ldAk20X6QQtWVgWSqWviO3Z8qmkbLdLVN8TgXosQF
Zjpz4ugk7jpoSlwLmUB/EXmDQg5E/6hv18DU03BCWTIfsNFI0JKUi31YKLCOoP1USbLwiJKpqNOL
kaXjjpvR6Fld7jnddf1OadGP5swKss0xlA8kM2YUboeggepLvQiVW9t7T3zX3CamYj4Z41lpM6tJ
NxtaOD4Ug1vLgb6Rn8wNPqwG5sY37QJFNenYsgZcrP7yYyHRvLSq0hXkMq9aSjJPZmjpCXbxpo5r
iSulb00gvkL5R/yewdxWegVgI7pk2vDL7TPzFlms7N+ac6qvlILnQbYxGRAJLUg6/vnGZnufH8re
EvMMUEv2GtiDe+5VEXizC208XHKdY5JIbRNgkrAXyJPwleCI/48car96kgqNdMn0LGEPdzbQeLxq
hYQa6rWHJaXJlVxwyvVcibSgREpKLw127NusPq8qmOgOAXxy/QCiPLpzyNcw5AalvxcSkuQtb+fr
bHx+ux2LiWqjoptum/FC8f+5WRQrfvmn2lxpyMHEIoGsH0CqbdA0qjR4zYRC7sC/SIq++UQzgmNS
6OEnnlcF+s19/GaoU238X6RpnBctA9BN09NXDH0MYdmb9AaEPoJu2yDaFrH6883a/TlkI6NakSZD
i2MQosCYvC7k944xWMVwhXqlWqE4PMTlpws+k+/c8pvh56NwmtE7z86VlSTR5CMlspdqjYKzgEj0
m7H0NILdiVWAPXwPIbj2nrw4wCvTpuwylCqyQ+kQvaqHf7L+vSwNCE+vTGA0iRLI0j1yhtKmkW6n
AYAz+k1nNcuWR/10dgeN6yEz3IMDVyN4ljMYqG4borkWAT4kLFzm3FTTNiDdrojv9sABtvN2zQ3X
ZLedRw51k+nkTFMJlX1zZACNXVa2LkMP+4/XzKzBbm9g1evym8IL2mdlBLTlea8WX+eTZ5M1Ns3Y
l6EWxfEfhk98mXLS/XuvdwApJE2y778t0hovq9yLThdJ/MQFvIJ3kjA4iWgvS6i0i9Euzvw+iP/y
oBJgOmtfoBUs/vgU78VTBoFiAP4RRVFulbLPcQ8RhtLu6dI+RbwhVo34C3E4Hr6m0f0HJagpbyLm
Xzn7Fvy2tlA0KsLzZsL++4uf4nSFaL5Znz+IIny6TbGSZbbsUPrDPtYZkrRQHk00KeHTXEGS72ut
lwlQl+O+oz/vvaHOMQc5XyeLdCMqh2KlESVpHBM+EIHxdSoP/4w+nosSgHBpvgkMI65yOzIqP9Lr
iXHt6iC1uAGa+iUXys5xZEoSznuLzl5gWhKXSM0ZFzTVZJSey3JvYTXeJlp3J5C20M9wxMVNj3Dk
FaoEFO7Y3Akb9FSo/H1hblKYbq5oNMclhdKze+dU2ubUK44Z1F4csyi8/uobgRY0yKyx/U2TyI1B
VwqMgo6yIhUIce7U+CWZOtbCVQIROXlMe8KT+msWH/b67ME83waR7Y2tR0wL6zY5SQ+SibuYsROf
UUeH964IrXI2d5ZtskfmBt+MNRhil7Tee5jRt0jrnBrK+asjYmTvyTCHNyYXTvZ9gezV9iGqhh+y
20BquW7brFZ1xx9z15OMRmNpMnOEPfUCqrd+JvMuBS8nkRicTPKTxezun4bdX3Fmuu1cl+Uy5bpx
mm+McJ2ePkVkmaLCQ7GnY+/0zfYIxrVzyYKK82g0TWB9IeC0dlVBbd8L/ACdbie9gmnebJHTt2aT
i7JzDSVUUs5srVQTgFl38C9DuOyHJa75Vr9Odzd8ffuzbr18ujero2RI707PO+vJhjVcyfd89X0/
v4c3CHCac6+PXzWdCGOvXopw+fc34d9ySgnz2EDdV9NdlA5Aj7pAX/YBxqVDQdTwZSJZ7BpmB4K0
LsYpYeeUuPqMlIjYvANl0gPzsZa7b0mm/OaLFCx5ujt2EuMMgoIBHHZRy1mp8W+maSEvld71b9dp
1pUlByKXlHbqmQxGSpZ3fFeqoNQIblOZkkX/p7Oc3PHiTf61PcPqWyPogOnVrN1tDvYT+ZI/WDWm
1HWm4La/iVm+buzJ0modV6VnujWSD3hy8zI/+bBBGBloO/LEyjmGwHCK2xzxf7mJQC5jsjSbFvtp
LlZEIylDlb3ujHx15zOc1eoBfKd4caFbU0UIFeXq9e1RqOOeBby8K/WJrnPNS9OtlXFSuegtzGwX
vB5K5WvtVC1plHOR+IRqCNF7ZIy2DK9zgJibhKcYdlyUWhg+D2jUfRY56pa8mk+KazTsW3yuYgCc
1UglryL9GIcPtxus6JAswNpJgM4byu8C/fcLaCAeZXe/mOhuxY05/nKV9yrGHFYsa3JRWroYmMkf
FF6B0mouFJQhQIOG6333hnGwrA9WmGmL9WyfD93WZt3Ww3UMbeWOcriHcvlWd2G5yc+yftgOu8Hm
3Yw6BS5LRMrro4CYxCnqjmb9uEByrIFvXSEuptASwjX/AzVq/PGRwyXpz6qf/+rFvVCmjtwt+urM
bioEsroej2bhKyammU9AP8VAqLw6a77r1bARLuMJYKXcbpo/a0llwHYIE6FpCDdDtEfWeeHWhs25
jfkdgfR6+CKx5GODqqSBYty4uhSTTDMLErqTL/YCZO0siagNZQPpYu94GZ136d3nzbs3V8swCN+h
SPxFWV1PpX1aQRXij9Iu3CxTgjJnTRBjJvvC+A8WG4K2Wpc9O3ChF73GyN2i4CFqw/s/Wprq2ax+
w9u5VncbiGj27qA3o1JVTcY2sLh8Ov8tudVJY7kaxT9JFD8wgxbQ7oh9IaQWzeYJFo3zdgc9XdVY
2cV8rB/sp8upW+wcIfLOhUJIEyKuEymQx669umQLP6jNNYhriMq6cJ1cNf90EdEVLTxJ9KOC2Ewc
0BICEX0KxnDr/NnjtzPvAM+y+j0j8KLf+MA7RUUkKgS4v4OHwjIOrNdLepU4Dads3ONNl7surDKg
D1CMTqO78BgZA3XXl+H14aOvZT8OrONYu7+dsLyjTCXCOKzQOcl8on6BUdGOj3igZNbHXUWx0Zdu
ZvteYNrhTYlju0ZkXNWRzpemkkhymZQWrcpGiMQfrmJpaTgUuUfTglHoD8ssg/8iKhCssw70dRs0
gqe/mNHF9eKCR1nQurmon+JJV3SPuDti6V5A9e7QxNkIWg2j1rhsNotz58qT5NGTXfWFErHix3vQ
2HoL0MAgtds5EdQzy9CYXMgFg4eD6waNq8hU0qkDQ9TjsvZmmaaZ+r2P8noInelI76eDx4Hx+6mX
9o0dQxn/voczYPuefH492PiDT4PEpYOdanCdbUtIhksLnSirKDSKnIy/J8lPMziPfuSqTPDSbs5Y
uwieFf0yXlzPEnz3LEvxWcBr7hfHBOUTFnqvMPY6t55P24yvqiq9YvW65btacH549y2oZoM1wOA3
NtQxNXaJOoxXQ/5jq2wpyBKIKRCUNF2n3i3i2mcpz31P5V7zKq8+axHUcO1HX/w+H1T9NQSzxAil
OSPW/ffXIg5GKkR9Jbg7NfCRqZQp/b7FoFUYeZNcglcsPmMNZkgMwViZW1qiyOleoIVyNAqUEV6x
bc/P48R4tJO3OMHVXewAmFEQWAJ4SqoHV54ChY8LyT9vgIur2DtbBP9JpFIDfZ5ikLKVSmLO7H7L
3yaJDjT21Kd5yk2MnIu4rBrWQ+8tuH4cWfv54DalXOaul9Q/lZJp89q+FfH8J113M+aiPwp506xU
n1n80M//EM5cN2YAoORun2qbYxl/mBpsWW1UmIP2aiCgiVsYPKLfMG+wyJLavDe1r2ae7f3Fnr2R
T283a21mM+hoPmQ5cr3OCaemE7o5W1p7GcWMC37RWbtqPINZ7sVVXrxD1OhwDCeCVyVNeMTsJl+G
nLbcRw24bgZYELJcvq5bnrpJA5CjvGYoX9EoWylKhEsUS7dWnwHsu9e7gvdfxa7694juUGNQpC5O
CvGioTtAvJHpijbzD1C7wRMeL+iK5WSlo4z+04KHhhAbTpGClStF1bEwOUikmGtCgQ98VzRp+rVu
P4Jp8kEvxJK4+u8XNjr6th4kBRsFp07ay+JojrMdx959qnbb/YEDCVE5NW9vp9qWjkul5YmnQrKX
BePXfwLoVAQFBDZAaEJGMUpWjKRosJXipViQNQZZ5lmENOUBQ5wWx7PJhochrEBUpchqKvJ//tyL
jGsFbgfPMk8TeNLGqBkUKtHu/L5lBDZYc0iNxk4PforzDsLEWO/iaEb3cjx5CxLSAfbuJtS99/fD
TpxXuzIrzJwdfS/0GYcJKMe661BNI76EwO0AMhAKGSqH9y5MDvzaVZSNp+df3vzUV0Zy32feM836
ksGcDkR02aQ7esYwW/djFBy8W6+Vb0u/sb+lIHBioB5YRyfAQnM+bcvi6J5r9ZAbems2qQBY9H1y
aWrdY1z67brcZJZJZC+wXLuJgQdhgh+QSQ6PQFPb3n3f/o+ilJ2tNOuet6Kji2++O6Yq3QdoQ/al
2ev/8Gg6aLkwQCZ8ujXJy4eLT7n2yRR+gJnnT6sZxmFCtNCzch1vozfJ+tugbPPmli7j2cFxnq4N
YqL90b9fOQ6H5eMi5VKSMcwPXTQowtdiPiqDqR7C7H5rtptsc/eWLMJ/ZOqS55TwCD8Sv1yWkMSf
k9jr2X7oYaH1A9Ylo2ihi0X5LKxPyNnUEdExUh17ixWqXZKAJFYbnDvZeYkpw7EMyrOClVbT+vl8
dMsalzQSRc07EOBLOZbSnV+gLi4V1fhDK85rWo1CVAVnlc42U/7+OqqbYCXgLp9/9YFRK1CavNd/
3Ng2qSs1NMmfrPfOCcEesGO1o+KYei3CdWCEuPR6xhA6QdAe5GGD/7MWe39fMfJSH/YDgfNs+PDw
gEKBCh34wNtH17z2SnkTPdfLOkLvt+RmRLz4olHgUVaEEm0s4Y2gT/kLrPSLkMo46fyYQDuq5GLp
DunvDo87WX6OaKof5RJXCYnk9kFnxd2/ZskJVRAHByCqPqkF5t3mnGhVYA6WUQozd3Yd1UNEceCv
b8UXfn8ql4S36xk4hslpjLv4VbykAccomkgZWg6GUDkboUZFdHZUQGiVn+sAZcJMvIOFbesfHXuF
grdi7abFaFQr57545EanPlZUGf/l08hydkpgEwOlm/NiK/byD3ubqCdake5n01kM/72tLdOfm9Sz
tjez+btBQyk6vA6OM2k5cKic3x8d26KH/sYYIBj0OrshRXX1IMbScQD+FUik3YLTZ21JYGDToCBx
bZP4lmQ4Qoep+sYHWgUgfTHO3OlKlnHXKsgFRkx1kSR02USEtH8lxLNTWdEPcFKfshWeRlrFSBE0
BUS/52EkUL8hWgz8K2XySLx3FfnXB3YJpzSN2wpFbmqBFEBgg0kifQ68TetKaSpS1Sbo97zb8ae6
b76ODgQPdzJpbWDr7S6sPqWyzcJkE8aFWFnespaHOJqru9ue1LagwbF7pkV7cAzd9BSKILJpZWmN
3YVR3pLyEXmjQYs67m4rRzr+qUV2T2DtgugKjk5WqojQ0DQHM/+OmHe4TOlrbty/ozGA8J35g2wG
Vnc+kc8DMwpeERBYXRCbYa4TY6ufsMYk+x2HlZx5+7BIGGQ2H4MPeVc8/6/kYkHXsuxEB9MQp8cL
4JAWFSsrzFcmwmUa9TzSZDhy/ryVTnn3yPaW0p9c72s0VqSayxEi1O/clQov6puWQ+lFynhGh5Hi
sCz45pZzQDcUBXLS4Krb0+b40c3JERX35iTPBCmigI4xfq6ajWo9si6aBf7mhRq3IYPHjQBW/Dtv
E3q5QZ3y1DkAmesnJ1usG9s6T4EX6lJT1Ol15W9WwTqTNNBobUuirJ3WVKcxGR9pT8yRpw4FrCuT
8svcqjjwls4EUjPw8yrXEdZg+osYnk1dDDsluGqpxw4AG9NREt9kSZ2pYJI4j3PlYi+93urz+cMQ
vkBgTUbVrHcdS5W3Uau1vt1nnxg3p14P0bk1h5IPIP3qHVlwjscGWD/gab4Rsi8EEiLanSjmkPDM
iKlHFQZiLCP8GxG9uKuM0L8JFUfabdjqjUw/3BhjMNSoT1sbhqvsFWHvI4vuglEjA7uXMmPTLTXp
1MdMl40cy5fK1gywSsZ1SzucjBAXiQopW4eIJwM2CKtPslEoTkGFtVeGKyRMagY9TBsx6xtGDYkb
ElgVgNrJl+nxbQxMdGTkl0i8RnCpYmTjzQS46tLLmG9ujYxffjA6hNbEkpBhh39adQa4GTk7By0z
0+KNHHc0kDrv43zDKIMX1MVjPILu1yY+ZkqLJFFyNG6AK4G0sq8W4iSb0bXei0pYBo2b4Y3MMsYb
PnPlQznqPnX76vdD/hWL03sw6AgHq5nr/2xurJ0jNP7+9Z3EIOIEei4wB9PFVpTZ8FoCrsARxL30
ePSAJq1QcZuj4u0OOzs3/7fN47Mkzj7gaHLZxoaMU7aXlT0TdbMnoUWegXaexuTAoo3rcWf2PJ1l
ivj2A3tcDfXRrsPZOZu65/EtawsbKDZhYWhMXwy5SrUJw3meMz8U/BQRRbVscHOwIyvno0M3GUiF
LlwEoBmqdzLwXMV8/yakmufcntcU/TuScIUJ6k7+bbpSIV0NNE4f1M/QDwAFP0/VQpiWLdt+apce
ffAwSgR7KJveQssAxl779FIrQixmiWIxb2+6oK5EvrRQsGjC/1uRzVIfzIfaOEfBcGLUMOawhHDm
s9JSoprClGhHGIIprcKRZFOwVh5mvaPQWshCfXDBH7/7WPI3I+274zp9WHML/nDMvYcRhuBXXoP6
Alle+7S4sofXQzT4BnjhwBBbRXtrWQX1M35QHCXQU2jwaqWwDqcYq9iOAWkGW7NyfnpykCBnjvrJ
5z+N85KhrXm5lUqNicAfK4TdGimtzcIJqqZ3B3PmI9YFwBXnUB2qdfM3Et730hspH42SUxyvq6N3
vlvXm58QZKj+ODVXo1ZyOE85PLTXW6prPypa8WBil7DUrbtYqZm0wTct4Yb8aQ5duTFB8vdCRRnG
EFh+6xUwAF7Dol+k2kPHRid+p43N1Cix/YqksR8zMngcc+mGUVFiTWICoTiM8YR8geRlAjL89crr
LL+I2OkukWaqbYuMt0hWi7JjHHlxju1T6zffTbIRe5YXOIopA91XsUkZ+Sd9578YyW0/oHDSYDi0
ZZFfU3TYcepgNB6+I6ribn4e5NwhjVYtPdfWTuLYYVzfSYCtnqRfR84SmRmyr7CxId2xJpvcVPQC
rt0SpExe/gpONYOOSijOW2AF0YLnAeZPBXzsKuerWY3p1uz+Vb3omptQOhmBoWMx1UNHue2bHr9Q
B+zthy6F+bkOiTHUNFfFyCRSbKl03336usISPWAqnXZ6Lgm03yALElqmUne1c0Pn8J42xvLRVWnF
3s/Zh9NmuaW0CF+LaUrVA1n91EsJhVAQgmb4vkCZ+DE5MfvVThhO+N/hP6Nz/m4MxEJXkA31a5l5
ardf7Y4GfrhwYFjjmSeZydJc6kEtBU7aGbUMmJfPFYuHLxMOhXQ1LzOjR0z+LLesI/gqUS7CqtNX
1TI6NwLrWOcwZaDAAnekYYEciZHi7Rv1XY7JNOGYMqIPGxsEuQe2EivZzzUDcODsTe4MfqXHUpFz
PrLaDL1ivbCVJm7BuVH8huD9D2njVSYJEdmSF1hgIrAehQ/IAawGYT+vwPo3gOYwDeiVPdC9ye1/
as6A6Va/fJwUwulOpWbTBENLQnHfPhBm5J9i1xRBaRwdQBWscJ6Ld67OwpcER2V834jNOhYCqV6i
4bPY1/N2RFT7WNk5sibjQlkgx4mGyifZh5GQj/l3xcLdGEvObJNwXCaPHu+c2+QKK5r49AhVpsib
ermJVpyQq3rr0tJta+OfI47lOEdnZtqV1fUOxSh3AyE7a0lSoPQnFdQ6MZUJIqNhAEgbEYy8yfMT
gSn/XFZ2Ud4Xbggn5DdP47Jwtl4VvXWs1Ri1VmEzV3gxKUyi/hYK2ShRn7EuvxBc29JK4PnzN19s
yeyYreOd4SMuZsVUXZs64OVvATAAAc5ApscGmedwdOESIu/HR5eDA22QyyXq9VjOOwGwyMDDv6CN
U63aJAXrtHWAFKc2O9v0bxlYP8MPeVcKxeagsjm44sws8nfELXe2OitCr/qiRn5CO6ciAqDCJdY5
InvXpBHl1C1e+ghRRNpmfPTy4ovgLLfzqUWH4jRhKmeEdN9P0LzZ+WDAjse4iKGm0CBJcZR3oEu4
g95mosI+JYN2Uw03KhjJyy7ZpGaIMHIBmppNI3nLxCy/qG9fyIoD82UfaxNgQ8vDTPeIjsZN2F2j
JoNvGGBI2gNsZsFzGxEn/2x5pxnPTIic5yDfMPFWG+UfEL+JOiYckJQ/ZdBZFLtRmiZIbM2iv/Uv
Gj82wzZKs5HonCHzaTZPTh8dHUNRjq8GdBmBi+u9zkEgvJZeE5uw0IHxc1Ty/t+Q2A+pYX6GbZ3u
/MEwLuweR/gkmPp2/bg9AVlIcrv6/wx0bhRzKJVu9s3AWbsas0lSu5+qKNOe/kqCq3uBlWpjyOml
+2z21/qg6cecdU1aLo3FfNEcQ1B0erLodJ3p5V+4AlZ2KO0XVjK/tDPvqqkPKWSfcQXzspzzvC7F
Vejcyu8egGTYzm4aefyZw/zCxPLk5gWfYfbqaATQmzSgxbaC8WOV9rxb7NoGOxvv5RAPRz3eEgdr
Vc6MzN5hTUN8YbAhPDKGBVNx3ae46za6H/M2kGcLYFzl62ojjZ8MC+nimcrhUAuW1grRAIwboRuT
RtrumRxb4VwIgG4ggXZZcHMISh8P/7AIVWWdPjPjWcZJQzGKs0g5AZcc2+MrUOVDOiYDRIS2/ZxJ
JKYtYanyAJ8stg1tBMbc5AyItA729v87UXFmzHwwuL5Q/XgN/nhJTA43cXKE8EsoYmoshbu6icRp
aRuSnCjDgeTPlEN78nX4Eutypye97iLztvEyWzM4UJBAaTYOIuvH1YryUuoXOA3jPNEVEoGAAw2s
by798zTqgiIpQHfOI5qndxOqsPAC4DyCdM5G/6bjAZsm91Yb7ZCigSoNeSZCZiUFSRSd7ojg0CtV
Cc+DqFzjS2cLevO3MtjtQwFznxHZVEDWNPjSQl5fv40W355gUTYoI7Vhb9E+9XY8khfdGfI46NgM
qqDMhNrul5GkDbU68rY3h+8VoxHkRaXUnCgnY/D0uYjBaiv4qzD01Ie/8lkcg0JVoFLAK7FUsGiX
tB57fNihTEUboQ+M9xiMCivoWY8L/txSe7QYkKDHEG1SgGSyLEo7FKgEWnMJ6OnBgM/GjWs3it7G
9uJbN9ynakZWPuGkt97MzLyXvQYxE3GquMlljQxnAFCPgZPZ6YUD3uXOdCJ3lqiPKxptQp6YB0AR
ukMTEx7jVplvVbDaDOHjYLp3PNTJYv56R0gDZeBJyYqUHXPrQLzkF2wPY6TJ7V2OUs9GBoVfClkp
iaX397gaJ3bxE45uELDVBFqBKGVJQ5LAV+ewhjobbzOWyvycPne3C5QBe1wVdGOl5VkGCcz6aATX
XzoVdYQTCTd8e+TsDbIsZOZXtnfwh2oemDkPC17S4cbAR/u2IucnGCxqhWxF1IvvLU++t0VEhfGf
PjUONEUTDwFUYF4Q4upfJ8Vn4BOXzj66E0pcsltMxz1U+12sLSdkc7cO7RuzO/Gfxp7p9xBNKC38
P7oF6OfIufwzk7IgH6HbKuQ7QMGlHIf+2CZRo6ihKw59BwJZQ0o0Z8zRUDWsYsEICfHPTRsNg6PP
+kyPPPd7WP97h5LqSR0IIcenmWnbzNVqqcSlU/036vTez45NULhSMWym/I2uFImI0luM+FgrDplT
x5KuuavVg1q4lJBZZnDI6+ImPJs5JX7zX3wmTYY/LECChICfvAAAeoIzXBhjx9VvpBu8G+SWq2hA
H3NEkgeDYRYXvq01Mc4gSNtiyDkHhnuCotgBI/qLXeQVno4jwx9jVERBX3YfHcqc8G0sC+JRaucf
+aJm97sxUdxVriGwnTZfY6WbhWJtwDAsQpWEAGposR+Z8FcJIsRsiZrNQbDSepFJkeUNvEOMOSIy
8db+OVAfRq4O+MNXgJK5UFjotkly+Eip+wNsDJj0EgzblfMDOAAhghxDoRthzDQ70imOCoBHsEVX
h5opkKVaq2aUhHOhE5SXbCAEedgJmQTtSSAAJWlF5uA2ta/imvCarWcD2rdpq9u9fHxaJNGGY0xS
5teEuO2Aec8KQvDXRfZTMsyz69pMh/3D2kNON7MuZVKRuu75yiK/YXbzUL4TPhPGp0pNO+BhW5CN
8yrSYXtGA9eXLgcrwsPCz82YFPVvvmrjfQMd0x6rWYnDtbzSSgrxzsrU/TuCpHtLdBHhEAOZ0N6I
UnR1aDmw6Xz17E1L141dNCd+1cFCEbsL7c6r+c47X7yvamKFRTzYuaF1kzlLdTEVKwZTN0TS57d1
6d/LowHFWLd+FGXKHYPuntfqCDG3Pm0msxRQwDbPzhEu7x7tEXfwdfzYHZiWz7cd0rVF7LS06zAV
KAezsBSFtzxYnVxx7Fufi6ui7e3dtcJOwvGy5xx+VAQ3r/TvAJtgCPxO+KwHbIiD6UhB1HCwlPkE
m7ikzJFWqm6lD53DkBwvWuFaHrJXx+L8RXpv5i5pCF32J5X3yt4FzZtNLQEkDSVRz8CzL7ZeoppQ
MXIkYScyyIUdF/oKEzoFd28eaxJeyiAeTS0QMA4Q0wd10i16eKHZjC3av6PC8jaJOnD5DO1Og6zw
6WH3ZWlagVuNRO6Q6oEhOOMA1wL404k5BQb6+iWfJF0rZCvKQUWOJ7gjp+Kp7J/Fr5UzrBAu9Qu9
Me+m5gAOgac1Xs+YOjBmSl14kcmQSbxazqE8f5qBgXGmsPdZHLfohEBF46z+682aMzFW5mm6YAAE
b/71o1TfT0XnaHM6myghzCSZ9lV89wSOc4hhCUlxaG4uGElYnseQDucarsAgGfb4q3bbksUaFVe5
l5u9aRR2KE5yxq8MWEyXaRc6b4YM8g2Yn+Kuhku0y+9JXhPuzk/QIaQqhYRQTYqtjAuFUEdmbhwb
4Kjut9y3qB4fPm5Kidh2T+hBZc6GSYmqAhq0pXs4jzTsUvg4BXFZWp0HoR7F1IdaV0xwIebCCZ8L
xhfWhScoYMMT1jahMKMFUXxfNSojxjDm5bEqxunUHyYvwlcVB7GF7M209Rm4LXf44zxfJIPT29VZ
7LdYOZTyb+Tm8QP717kfT3zWmFmcfLHwW+tVGwhMmKQQtOwnNuIk/3dARqNCBLBrZ1HgVCFeoOfH
kAgu1xHthgBO8oT+51qqOo8N+lahaw8NB401Eo4Yl71CHw5FzvKYWYgxsdkQ0yiA3vs6STNNhwun
8MafY5dmBFbJFNIKZzMb8Z8x0IFfcXxIakXFB280NMpxhHrdkg1VbAH9M/s/4wGW4SC7D2YkdcmL
ooeDnw1wrlUKdtq/9PTJM23JY2P4Xt/HJ1bOV+U8D5QYDKvqNGqIoZrTrZfP/q2g4S6wQ8UAOkqp
E/rWwPLX8i4ZypmYyKij0DGidwvnxiny5AISjLKHNakUjNSlsb4tq0YjyiagA8xX/+zJBwUs4bUK
p5XutVCrpMOoAFRDI3leMuzOmt6LS/K2hrBzLBSS8uZr7ZNkqvbxbNJ6I+satbqppVJd6BSScidu
vGsHwR4aSytHe/bFWzT9BPKXxf1RJg8URe9fU+mRhEfZPamAfAQ1guij9ORmedT1x0dqUzkhRYpY
BiFf+s0jc1j3i+9LcIp8CWyhDOqGjyBK+ONSyO/BNbGCQ57NTu4Tl0NciAgBNR7LJMSTYFdpVBJA
bRIDnMNs1B4ziBflP0WjXKwI10FJ0JGsCAY/jOPIG+SXBvYiH8bnLw5TCVqZ9tmJADk6Q74S4ahV
rEyBvFqnw4JOVTS8+FDqWFIw8ul0+KmH6laJ+rKQZ7cPhBY5YC2ephPpe9IdOQRcOVtVYw65M4iv
dpW0GwfkiNlXPrnhYFYFCgovYio/gwk+JLM2rF4Skn8XyUSuhiPJULXPayujF8LLNQ61jgd/klXM
WTcGBuVwG0PtRZ7XS620RXkxnmlTApvFm9Fq8fNMoTS+BX5b/GZHvTdoJxP7d2+HZUOxdMBnOTau
rltGzTf/D7sJ1vd3zaconuGvmPNVEATCTntkBAAxIQNHh6rG4hd7YLiYefUdLmEbbkQdJMBlZ7h7
lR39UXcR2c/dnGw1fj+On+S9irGzAvodnO/Kv8U/BKsCooyLVqHwTsppZHX2czCJDP2FUXKLUDNa
01EGX0Cz0z7+2xVVSOQ7jfV8WJLYqAD3VHlXK8xbmwulNcszx8ycsdamjrqA/vSAcNhJQvQpPJLW
tytf5zNtZ5jExsQ2PC19bTmmwrFEdUIDOttS6vu3gqfFZ+lfmgxdkva7JmfIlGhDZBpOstpwWWmx
G7sIR2gOFy3QH6bmwo32MtqE/0BvKZFBp7cHem1lYoOAZz+nHjk2KaxAgnb8pcMijjmaMKIB66zQ
z659GNNZWC5986dFdhKBNSjkn3eT8XCIsnZkuJfSHzkD/oZUCkWeJ7VK/k8+15uR9pOjU02D5J+S
uMWYtzT9I64QUtEwROOgqAsFfVxkGfxUNN0Sl0Ynaf+kOh82n4Pts+r93HcxepBqEukk7ubi3OST
hNiBCFbw5Be/Cem7MpAjPbgwTePOjxuoq1EQupp6tJRfzRFH5NcuuHmAFlcmSjr3RqJ53QZ2EGsb
T0spNuzDzE9II78DJQLilas+AfEIfs1mR+pa2s7vfTMXfxdGK9dBo6ZJZ6SCGSnP/+6TWpYUE+Mv
Drfvd07Led/uhwrKeS+p3a5YxzccYemUHFniYQEWOsQzDUDUilZ2Ryaz+sn2uugmRJTBUvu/fuDw
bhWFpUmZD3JOsow77Nzkr67KIQ0GoGwodkJLgycuzKOlA0YkeXJxa0Xf1FMVFHOHe4KdbB851LDr
ahWzVGG28BhdxhDen96fHbXsB+FwMEi+DtNgEPJyx65i242FMTHP3TpnoxmgjjTt3GyYwsa9G82A
Vd+Wn3Wg1u6cS2+ggCL9GdFKvsQ0WAHKl06tmYwWN1kO0QoT7PLjoyYy6DsIhHiSwzdLJKLpMegS
ZEEly48wkQ6FT+dAOhSEHiJE7PGXH5ERnl1b2ngL29WHnMrs7d6iIDvVfYWTCJSv9rec8eqtCWg2
rY4ak+q24XXK6EGpTROX59ncelwFGtzn3txROkTeD+N3ycg76m3zy5o+zfdMio/atGsSwwNY2MhZ
YGqrzTL/aUpKIqlbeZrkfhcI4jeqDeAJxBbo2xZQN10uNZpOpn3kD2igvXbfJj1Fu7UNFDGDWTxk
5ONKoMgyiqa/LaQG7M4JTeZDQzTH72UAxHGBFWcLRIdVaKl6gXYad/XBztSRgRPgzama12pTj1kf
Jdak5YmCQsN2jlYIVSLXwiWd32JnGeOMqZkUEPJCzskN60p0T+dUWUeMhlnmwX2ikEBVygfJkg6g
gsJWqiQ1ritTfQDZbo4GYHOYPQTkb1qTLXl9CbXM3zNW/9CnkLH8Wry8+0xWeHV3X0iQX7pIt7PH
ZXFaz+ek7lIzPN+Dh49bfV2flqlDi3rLO821uegXBHfzA6VW+bojT80J3GPZ6bc6Z8suC3WrKRcJ
yz3ArCmddWF7fyU+OBj4Voc1ok0UBRtdq0EcIfBfXUWHS268D9tc+WY566m7IFVzgy6jP8ONJZ8v
f1Cbiq84+fkbxHZUFfnWq55njyh+peax+lg9XwwSZAhLEBMKP7AJ5vpAK90LwFsT6u3o14kd2wfH
IKhwWBJwfMLnYGNnvYd2E1EODPgFgToas4RsTMZMoGzwyckK1QK8mlJkvJ8KtyHvuF51YYmDxZuX
YkNzayhCb7OWdoDiZ8u65C4Ag4/jKxFe7qfKDRY86sIXF47StVEd/CnBWnzlQkcf3zwpZlbi8hOC
USFA12Zsq2L7/it2p92A91rURoi9qBbNSBSsQ/NoGXz3ipyrK++ft8ei+vj5lPRvBDbO0VhUmRX2
YhlJVC4ykJYzjytOumrCCmgelwU0CXFI7u/PiovP7ciEbtn6rSiWyGbMu+EJdycmj6sVc9qBxAt4
6VdAezP+ib2JbDZgh5R4702BB1breQk5PstDBVN0jtz+61LNLy4QEXTZekQNW8HhI7YGw8ofRmsv
keFpbAqYF+jcH4D0VRqWKTEDKOZywErvgUhzcVkvFBeyP+7FQVU6gJunzZpwDop2UCFP+IPPDGgT
aBSZAl58tyrr1ByTzHsK+9IFTFuyEIkjumeY4/UjxZ41dUTmKXT5fdLWVYegomNhSsTfbDuqxlfc
Q8XIcWTc715HgWCBClVu3PrvG7YT0N56CXkhEcerZR5FbNw30zjLxaC7eSoUfJ2wckGcv+iZDPMd
g6TcD/6+6J2kObyk1yde0gGwiA907DdamK2zDg+C7YjLl/6m1s+XUFoMAnHi7NMCJoMmrvIqGsSb
N4sWguXAbEz1/uGcR9G/CjMkeylpV+MDYIIQfZHWW8MEgBJkLC7hbOMOmZmzllLtFTuTGBN5AW9L
meWgMfPX1kXxDWAPBZiTqUgITCZTV5xjpLK4jMcs/qyLCD0dso8gvkShDXlsF43duG3MC5vJDKuY
x8fOgqPcENeW4HboSAP+JqI3vO8FvDhumGsfZ/aC+mJxWWQmapICe+wm11BVgE0UOH2AGqDTZfLk
9G7+1d5NeZg/8HzEEPi/J46pUoeNyjoLS2pnYN0xxr3XNkifvNiOA7oy6iRD3S/n8+bcq9Jn1p1w
uDI09wir/bSfQ3EukF0O87D20RVk3lcjnpGajP5D1OtU5P2TUcZL8vwHLpUN9qwmmf06bClS2xEi
awCDXfByLQ1o8XQnQ8uTAtLFHE5PxdBEli2IYuz0t7l7rO3ucPab5tD9g4jGPRlra0cUj3Voo311
R+fxpaP3nNDg0DhuOTf7fDUVlP24gh3nEZeGdLMz868Jn1n1JDEqygBDWBPUfJ9/H5kxorTH90cL
Ps1kpZY4JaMf66Vwd4NiwDL/W1nijz7y5UVqvzkNP3Kjl/6nlwdzY+GvxEM8eXN6/vUmSLcD+90Z
kg+C6Kh98i6VSuk92EbYri6lArc83Y+eRS3kHraQE/p31WKcFmp7ZQFwjeVV9jWaVYPp8yQbIz5w
o0SqDMRrhXf3ykNgrgRa9ONy5tkKmeF+IFkj9x/Rvh2BqAM0/UIZGwp3I0LCyIuHWlGzhPOnwCTV
5d834dhyMOl3S/573ZQZlcHb4SaDavwMh1C12clkz4SRUoT8UfPlOn8u3TBmk++lEVqmtpq8wen7
jon4qZ2wwRSsKQs+ZjrEv9cT/6PMqcyVqOUbvQqDCQGsc4e55fALSGmXO5sFlwGO62Ip/Vc/7bfJ
yyX/m5g6/bQpk+6zOlJNl5a11jMwX962G06nX663+cELUSHyc3a98iecUINtT344h6NVx3H/qZHZ
N3rBXKFABcA1rgOlWuWfJ9MqqOyecBDiP9g71ptJAxEXnEgskCwziuNGx52YZaNwmIIlJF3thnvC
Sy/k/VFwp+M/w3GsBbmnntnD643RCkcjqwF8Sr8wUh5WPzIMfQkCM8DlxunF1cxQAiHO1klU702h
RkNX/KeqObRBfVQxV6arqgvQOfCuXH6sOw5XIPTH3sxfT9X+8UjqCwSH9H9/w6vyZUjQdMvM0znc
E65vXey8TeacFU0dZP2Yafkee63TQhOQcvx3BEixfHPohg+Ew/8tyYl36V1/YglEc9ST2FhiMcuf
RdVoQYRZxEe7JCfFEEkKaRqpnTRl8xLKZ4CXq/1jlh2toAGFho9IPeetfrB3m/KvpOPRe9CtGBFr
Ukyd/JXGe2+r+zTFz8b8hL4b14g9T3IIq4D7tmBn5qDo+kafc8XoAfDpGhjKMXfKZD+kXqN4F/Fz
n9QsuOcATuhJWog7lzUmY4sLj1I/Jo7QSd2riaTDFSCEOsE7CIjGI5AgEcgm/vhW+2vzSmkb2eWm
UpOIIp7ycVmtJxFIWOEHDX1+Kj+RT97+HRONDUbIo4e5GwcZKwcYPkjHx6WHm/7TdCwBaIJQ69ew
+GlYwQfITdOignwofqsykTnYuY9BzPhSn2+ULru74xVJGoZyhVRhI/wjLdIryuKGK50SSjF53NcY
vKPfS80UjVlGv2jKY4UzeudnyIg0NMcl/bS1s+rM8subocHZD9v7EtdaaFbJmdfNISfpGqC4N24A
6MFudILA1nHyu9g+HS8SM4T4zqxZqJGOboJ8rdTQzrePrjYB3K6Odt0zehtGUicXHMB8qREk+fQ1
97A1OhMSGQz90wvaY/ywIq0gaES2rF3Ei+SkL7622xYZzSxiH5D1+qzEL7CLnLejELDKCNapPyf6
yqRzPLJp3tCm1gMSxMGNbrVb5Pew3YBQndHSOaVTQQAtHQjQ4uxD1V/nUS2Ihln5ig7gwmQZ6a1U
HwQ3gWtrHGcQT/JauRSYa6b4QypBCdwN1cuqyrKL2Prq5Ree+PDKRwWDCCc7PmNEly58+82zeZAR
jkD5IcxkMn44oFYgLGNYP7YlD2/kZ208J0Qw+D/Ovflp6vDWJww+ExPC/0NDtZ8IMP+bIq7rndv3
CfQRv2PqiLDmFsTGjfBpYxVXU+vzb52ODXEEeFZZBaWbulpy47scVcfskugjtmx9e5jkE068Mar7
086i7GMKGDDZaYwLKZK04LeCj+oNvrlgQHzLzWq4LsS2FKKRmSTHBqeVgEwlKnw5xUC8qi5UmqSV
OMvvWVPKiyZx/L4IFBruBKc63h1EbFbG+/FbIyNDNWJJyJUuHo5CBgdcfyNX7q+uouyZqxriZs6F
voyAbHflrmvRoH+URVFj3+HDZ33stvt1/TzpLCGpKccUReKpP3oqnuFXyVGbzCWmxQxlaXaVmvwA
W5r6Tr7Iqsx/pr2PkaGQAGTauzTMyt+dodydsa1QfvYSdUy0y1JelysaCq01qcW/UBbxhpmwR69I
uvzGW6QKZHVzJ9XALy8nbpOIyJmgUlMZXUU+nWpAwJkzxCe7ddbGafWTjr8Zl1oGo+ZcOzZiik73
rdkCMuPRI2ctREyTXVEddlLmeUCffeLF+1tlGuDlECrR92aGNVxAv7Ansz5OZa4tz9eKfxtKNrxt
hzo/+59OEmL2WlYVEOoH0nedUCk80THqo8rYJGXbtFEB6otAQM8wIe2fVBH7/nI6IVPZ5L7KKNBe
mlPaQfQDBhl+YV/cOS0KDX3rAfXfmPtFm1mQiZwIyDbDhJdTl/x49dC2RewO4f6cdqfLuJN39uCa
YV4nw8dGakpQYlpjH0XnZxu6fIwmbcYUMfUkyvDbvboqJQdrd32lgtYBl34O/mmR68rsEBsKWvP1
5CiZ9cisyEA3oVBbtA8yGvetCn8uJUjc/hsajyNKgsrcWaEy3hMI3owaGDKU1TI7a1hpTp3hITK5
eShmDWdN6K705tsNdIleDoPJ/z++0sOJCI1bZ7TlN2UJCroPcVU2w7D46x71vv4UOuJ4BBx68nGA
k2nmEg5733lKlJwUBM4QHHShyHxgLgFAMjeqDZF+uoHaKS2JPi4G4lDTHpG1V/oy4c8HQb/zt6uj
5qW9JW/qC2lHP4lj5PbCgDAgPywbrLQPoxL7R6+TpV6W0krUJ5b/JzsX+PMMOPj+R82v9nEGCGQf
v2pcPctjMJmxR2HLEl1eqfr712t3oRitGeH8a0wpX3vbzG5S/rg2aTW29yKtE4+PoBwWXpCgz27I
ODrK4G7ObJbAXDQTUFod2Y6dzUrYPt+qhq3p7jPrBaSZkCoJtpOnkRpp6RUZWQV4OJNPitPO83mG
mFZ6u2aalE3omW2FY6OFMLW6c6t6U+AaBh43U9aRfUcDe6n+FWf00qh+j1mcwyLz586GRqBf0UlO
Vw66v7eH1rgvMsXuBYQeMwvbtHlV/W0ESli+Gl8mEq1+9C9wJ/5co6hPo9RpK+mcBfrAp3zvtwlP
wS3vlXUem3X9jywdeGUVwXU2es4LRWESPOXSMHKFlJzvHGwsrv1FqOS5Gof2iAN/A11lu/uhcXoh
QoHLyI5RF5FSCP7mMsvuY31IacUtl0TyBUh9/NuBzXDMVORNwzcSy3Ue2nSqB/wkph0orekm3HCB
5Em0xtVXTQD8Y6S67X90drSwEFgJWkwNeL9FoYl91r6QlH0CBSXT2iyLMF2ecHpgZgwrT8wvdKf5
w3V/AtdYMXxK+5vjV/2s3d/oWgRhb/dULg2LF0urJ3kYUGnxmeamT3sup3JD1eyHtGIBoo+z4hpT
UvFDsvTAYAdLtQej6l0OPGVn4RXoSIZb5wVUXw02XBwKBj9NEzOkmrxdR5qQnXoq+8m2UdkNpHcJ
bsn6vGfPG44SpoXz5osu+rHS6GaQC0GyW9Xr74irRqpNtqhoe+v8Q0L30o+ImoMMuuD4bsKpN2xD
0JIe8ho2+t+xwaGm80m+UsRLSLPSBo4FAFIp2ioFMRyEAY5FH8IoQnMfqTUqmVQZcvBqfdrFxPyx
J6V2H+Ovuq77AEKP6BKhpZ8e2pvuOs0XIdc752r62vOCDU+ZV2YlnJeHUWbwtKlDYA2u2fsQUUSz
EpoNmAFhhbAHH/e+NYhvjWhhnTSXscgjMAj8+0rdNgKq+VCtQuWGRn8z5of3rMcXrDnMu/3wE1jH
gwFA11qnTW1DEJkrsfYpvMmUq6nNEjUtlQJ6O9s9gvDIkCJ6wZqhFUG5DGbjb/ikC/uldnvTsaVM
5WVcVAjTUGHiS1aP4Vk3l2TNfwX/isM32611kITnD4rT8MiCn41oZ643BI4ykrdCXP1g9Q5hJaW2
u26ACZqrlQZW0pY6VTepUF4ydctLYf4Km+o/36N3rI3sXzIJpRx3dabE1fx/bTjZXzPrmetR8LEZ
WkwjmPARwrmscSHbpzU1dG4rl1R7ae6Iu/rH+jb67Rx206dEnacIbmeFNzlOd3jgGeJzGrGj8E5w
jFIcH2YNzi/JnfVbJTuXK5Wu3erVQfcnIS71LIRtNnqz0/wzrtrRpg7v2dXO8R7xsAHfYHU1i/pM
BPk3rbJrvgagr/Kq5+7kmEFynO2tV3wDRtE7dVG1hOvsj+ji7RtSzdbKysdaBDJ5KWe1tWoaC4Ab
RVuIr7H5UWbYLfg6jW/b6w5S0t59L0fNKIdmlVevxRbCY3ge8wgyK1jA9IvIVmusGbshNZHUAkYd
0R6VHCF/+RpGeYe8hJ5ZpJLHmO5//dG7yBcWiTjfwh67yBzX/6JaoT92fdTh/pKcSjcuEOrntVnP
OhyOKORsBSiorDrnocw/0WH5ytgabOp+mDXt8rFSyEB1NeTZnwHxVKphMhTbiecBKtMuZ2a3n4tm
EPoDT8M+dN6w6iqzSakUQ7IcWNvKBcLwcBHpKNkR1LYvjexTZehL27IvJgC52fYLXgLGFlc+gqBT
rSQy7l1G0iAv6rIEDA6WTc0cpYfeEROH3SIJP624VMCJXCV1T/IA26E/92/3NNBFLri7r2C3Z8b3
HWx7F21k5SLVcdOR35QcA1pQYyPlf+1+F2tjbQVAnUTf89xIAJg2cYIZCRq2syiCKRg8L2nOPuOV
ugCncp/ukYu/pI/5OcXJdI+mBy/q3V0Vfr1vw/YfCf5t6ykkATbslfB8kotUY/DeC+zFgZ1nnc1r
9cc5klfb6ZUWaRQdRfIUHekbL77Yd+yJnjxH+J2tDtv0H0S0hy+qz+Fdv8+I4tFo6qe3bUCW6yXo
UtsRff20M2MECC+16H/WxB5n87KhRO4immsS1jGLgAVOjKA6HbGoXieOiMlh1bV1S6hjgOrr3lnr
zvubFJ9She7fOHli2OnZ59b4HbxCCZJl34AYNjULdvArA4qEJrU0C05NSlVnKp1YFifQk3OSwr7l
PNrEWM6ds9QBbHWpuU33X2TU9IWubI1IO/aJvGLBBY8rc8MKA+mTIDQyl+4oCUsCMcss5+wwZyWY
U7DIclT2EYv4OmY9z9qpyJd1cqSOReMHtyDBOnXpMbIdACxPa3KTkgTFlxAgu2m0fHa6nUh1FQH5
F7vdkh0O5sXjJXeVnLVrARfv1gmgkp1xUiMZI604buBOnxPzM8raUCdbtS6GHpUmG0oJK9K2J7pW
/W+qaEyEFcQQ1iJan/Umj28bDdfxnv2xN/xX1JnA+BXk4MEx7NPfJsl+MlerTftyMBt7+TEBMEls
buZ+iQLq60i9B8tNsc6Amt5ZgXFW4JiKU5NQ4Rgb01mqr8Tz9kuRhvND8GkUhuLlxm5B1XVnMDPI
uyilc7+VXqMwMPaG/laAH2Wkx1gprlkAKliqyW8/ACerLGUm8aeJXy7GtF1VB57o+FvSvJABrSCE
cT8vw/SnTom7ASf4XpBguSp/KG93vv4FQBZ8Lx3M7Cvmub5BMmEtt1m0U3AYWBC6705kYeJhChEL
EyOzOpUxhaC18wcIcmo/13+g5idnlanhr9E22glf09Rie5HvK5wJFRX4Yw1EDaEu42nY/Qlvenfc
kfkoV0ohSCG2PefDTh7IUNX3ZP5N6fTCe0OBxd+Io/ZvtBW6R2m/J+flPXvq+SvpR4+H5inhSt0s
Yuf10PBzQxbQVhd5U+N/LQsqTtBPqbuS19WMz4AU5FZzgzKXEZ7WfMdRFAMsjrw43/voELU+tGbJ
6LUKTaSJzjmATFoLxT1RYko+nD4AxjXvrn3KVf/k4DpBo7Oo/5wx/6T3Xb+gegDj8kaSZiVLNziQ
BvM2eAL8XUpv31eOiqwVIFEvQzFA4MSwEcpMu9+d2LTlOkvSyejyIsPuijM/Jd0Rzg2phr4RDd6g
p7zW/1fQLKx74AxHSBfI9wXhyv+7uAKFU7bCw9CzXksOE8cql+nmS6HuDeYwKTHBDTv/56qjiZce
jXX6Ps8XhMeR0pS/yFQEwdhYIgWCJ8lTsaoTwHgECPwdxTFu/35DmjtWhWaSWIFNmYqVMeW8PT5G
6xnNOSewai+Xu8g8ZDGsPra7wYQ2Qcp1Q45oK6WW5PGUd6dbqNRtteE1PRSnzUZZknJzAvP1Kvlr
ncIISaXDGXqv4B5GbA2yeq+bS8ExH1haCZ4HGek5BvcDjNs0pXMoIdC/OnMGS6YYkhPcniVf4Y3/
Rdw2/erEclFCKUAeZH7kSuIesmd6BrykAyAhYL4jruuMwJR3p0Pvg27m/lx+pB8yAT0sUCbszS2H
apJXuqXKCio1Blhme/uDoOYkQJQv7iQ39wIwT0Q5k8zF9Cc62hq+/OCd5PN6kQqO/pWIhAUZpfXI
0T7rtffPGpF4xapcpDm2yBa7gRdmaXEppb86IhoasyWdKU6TF6QjVr67hAE8WELjupv7M7BZd28U
qFNofLrReLSrFHhnmKjdsfgJNMcl8v0yItJr/iNPs3978doIQJVA1vMmwLuzMVYVY/mf6frfQduP
aKhriCE0+S3gDilQBsI8zdR2k4th/tStiVvVwalxbjwtl/YWvXmXDTPSREUOUgT4h/UrjNpaOrdg
xFMkk0fui6w66ObdvBH0ulRm/KDzIa+x+XE2ZZiuep4pL4+9YjkDedfI5OY1B33uERGqsOLY/pni
gtue5WR+sC1AbOyBa83h0ljDL05GST+l163hEOv+EwuvHQoeNV6/AKUCDBUC4+7L5IzsrZuN6dxK
EwX0dPkHmEOi4NZNPXums8Cbq9R/a989/W6DcMUlAIByGiK5xXDx2Hk9IEDl5Qm6ZtJVruJYfrnn
NGz1asYG3XrXcvok5nI1TREv5Esl9vUkYPZHCAtG8pMqx5wW5tddcY7KkRbWGaM2RlJ1LrPGijeH
GBOx05Gb3eUGKyEelN1D5ubunAxYdBfvEyAICH/IAmHUCVyt9i4uo9yA+4WJmxwajOIwgDqRfg4B
FXhYnXlM3BpgHO+6d2GftWS1OkIeOVSe1ceSqMGJ/m1SDFNj7w6ZfHxBXjgabsyt4i6ylo8+5ges
mo6yVEQaG7WuSHOWhzplaNU8Z4sZx68FFsNEGiPnlSE6SJxIo5/IBtQL6ZTEmPtuybqbEA6unC1b
sgNdymHwPX86aaIcwQ0SNw8wH+DqlktbIfyoKZ+BoDY/UTa6QfFDSV2KNnxdhdwaqqV52k9IbUem
U9A3bbV6Q7Xyu6vUTLUVYwvVnqXAYiE+tSenFGqcfCnmOHwZKasvPrHCMSbXxQ52TDLad+8ZG8G1
bx8ZKT1aGWR1wB4sVwQAgQDZ4/5EWWbM22RfuhccHq0RwbWYZgZFHh0aQ7qYoEPCH+xwHhvuxbsb
nQKyUe3QkvyMVY20BJlgqMy7pmCNBc0ycywDxgfctDhjL6VRJJgCc9ZaLbK3JaOSh2TUtnClf71s
BgnzZs2UP5nMA1LKrMVMBYeTJY3BimoOySUWxX/WEoYjL0XwzOOkEBrik4HDCSRZFwa79ZQcbYXC
119/8ZlL6eNlcIfZJFEuueFqGGYUXDOpjPR7eK+DRQvn6QQ2ofxUwIOYoQWaeL3QgvurpjHlop0m
BFcOPULhf7B1AbS3Q2lPPwILO2G0I0Ivj8LBTc7Iuorn5p5x/Zr5fdcSppseRuz2vcCpy9hj+lnU
H5AdU/zrzdWEJeQSC2g3ItOB9If3J6nle90sbCW+nFL080LLXRE7dev+UqGllFiG51ktPGJqVBSW
F5rsJKzZmLeNKQ9wQRVAHSDwlEs76uuoOJ8Lzdf8/vrgFqhC5dQxS7ouzTl9uVKEfYCNzVHy604x
m6nd+C+6RxE5L1cWpyPnttyBZn9/mO2K7hgTXgxntKxu2i5ol0ZDd1VIj7s1Vh4QZ3HvQkdKccql
hz2SWBxhVm9XDu1Xbwb3LiZLnIqQBMZLgdjITKtCqkgagEKpziyfENyOhU6r1c21cyP7VyHRDaCA
TLD+SwBkmrl7ZCC9uk9r9DieOf8oQH3uYnAREdAxPc/K/iUKyRAaoNAIhqKjV0IToq0R6wWmbSZE
sliHkZniBXbG8rb+Fufdqfgf5Rp7a1bouo/HkBiRoO/GNsTF6VmgeSgv1LEoaCaYAX342AqF1fWB
IUyTs6EHrKPjeS9C49+wSzZ59I9WaSqinzg/H5z2+DTAtaDLCE/Y3sFFZkOt8ccZpZniNqVE4P9x
GpC0RFHQEgiLe/up8UyxJSzo86ILtxzXp3XSlsifXJpodA4YGXgbQdVReAhaZiQ9cqbsawW0g5PM
cWQw5/i813wkTrTTfWqGXVF7EU8DtVvs90d7GkEp5dxNnvUM8rR1ZVNoDZTuekyAzDbr1HUJC+oB
70EIrCGgvcOvpT1L+EOIK3o8rKEcTSwoI1SwN1I5lxC5/MBivzWmwVvFdRrBMA3go9IsSr7rKWZZ
oYt6MbT2Wt6HkKyX+Jtxn9msxu5uM/96XsF759o8qD1CRpmJpbP4qPmB1sxWv3HwO8f6SP+Bnfzg
30u6iQs0khk0b7dQBYNdWSKymyYxUXP1iWqQVufe3I4gUbpLvjpnpPbNXMdaLL5I/QhrPbplxMj1
Judzlbfe7PR/zWUvC2xewVoGcpLFAHV36v+lDgzUHvO0dP+liD2JkOn1jQda5+O8xqmPdEnhhp78
dhlhKCql6KZpe0bihxYJOSfUrzcNMuW4pLNDIufmjbazZzRjKX9V80512athzKT2ckS04K6H6cFc
V847FSm2gNFOWFjzLoYwn1qoipwycEP9AMNOSFS+XaFlOmLryU4Y6worU9XYTHBEEAHhmaMBiQFh
y9zTQDD/c+xNiahrjYuZmWEU1ud7c25piiXH/4MrhpPV4qxw1uC+KndVX0XFEfEePa6vZHJoUo/r
PLc8DfNrm81WrL8V2s+ZH8IcwAQOXc0GfUR7/1ZnWA8iv4OSj0GMQLfJk268k+uXXy4+Kk4a6eBL
8G5RPHUDSJpg9dSlmVhoSmYr0i9pXtI0FNDn4r2tTuabS3o3mzfZNZdAodTxSdCiOMU9LnwPScvw
Q5XKdAIUk8H0s4dFxvV4JcSGN2wzL9rTdawGH/RFxpLnb6BdVQC5+tn8tSWdc7r3bym7CoPFKWBq
QZjuC8nBk/ajYpY7heHcoiHX19H5l+Sn4jBJCjpKQAP/p0rI+3Qb8mRERxnNfRB9ubI48snxRAz2
dJ3tLj7mRQPbwpVe1RF+q/GVVJtUPNPj62qftXZmja9SIQOufMGSq5mGiqfH89O/3pB+1zILgKGD
kkLIIYDZk94glGpQT0L3LT6g0g94pCg4RGB6tXEpR4g26/ENVTFbvSHMh/qRA8t/OL1yDuF56C96
VMn4y+ATm0yhorGsIWRHbOGZVkb3bWjcsy4MYgo0tfUIa15trxStoxeBu2rRW/KuiQ9CD03K/Zmk
UBjZOLqBoMIh/Zpim/kYZdJaTQELvDwhO13d9YNqlf9yz++5I4qvoJQdLXSECzVNiLFbFQ+RhnAC
7+bAA1F+CbUIBoc/sx7RwTFZrhT5SkKvC4WjQR9vbLH9ZTEuD4fSveLpL0jmhdFzynF4J9TyKDZu
yNeG4A+bP/e7PjtW+c4mDdQ8jNnALVq/zXuAJvuxysnd7uY3Adi1DxS0CRnGwc+urNvdRfbJv+OJ
3FLHgRQC5iDhY72VE6l0rdieYONcQsnGcSlnO4WOqgWxb2FfDVVzA1XX1VgqxfXYGoqa4PiqgAJF
TQKFL5zu09TaqnzFAitftHBGanzz2O4VU5+MjH4oXCt3Oshic/uMhVejIO37F6pSG9puUVTsJi0A
LFzD4pe+WezSWaKHocjFeuB2mct4sjsgidJWw+AikGjJeQK3C0B1V75h9t4Qokp1C9JCZehhFo9C
bgOXgHNXUmLiHZcETF9geOUXS74+tcetkvWxEuXRfw51NYXY+XQd8UgKKn4T6lN1EwbD0QWP069/
foBqgH9A5JjKqS2CTJe8berwPO216GnkN5ro0rp3nqTG5D0eeFKl++/kjLVc2BMk0YQgezeKwqNS
ywkB90UGnv+YV06uC1LaL3MdccSLnD5Vh0KWxfyq7C+F1ypglVTyJKxUn12ANH0TEGp/POSg+/ig
Gleb6sHKljD+tQ997MCgwU7jt+z76qh2+ET6Caeb5jUAXKbp3CdVCdxMIFt6AFagcbYmqq+nimyM
VdfAmKmjdrFG5znGj57z4FMo1/17i3zUsBvY8MEe5GzDq79H0GWmWCAu0ZjqpDJVsFdUwgyL7y19
2wECp/4GNuO0xM6gQyUclvwEgmvW+Qlnz6h0yNguLcOeyBw8DDSpQb8wXX4UAXU1R2Rq781IxdBY
JyirxcRJOEIH2Sq2HwfPSXQSVZX5n14+cUgpSM9gqrVImk+ooDoh5Xtzk2xxzkncV70zMlj9cS17
WdsQBX8P7quH/93WPgWGgS72yGPSbUZfxvE3jyC4XJ3SIsLWYv3HRd48OlN6dU0ZgJo5dKORUC0r
10iPPxEL5cFwQc5CKc5hyBkrbOLUDBfkP871L2BXeB2/klOWBHM9LgjTLCZUJw+Yz9sy1W7ghZS6
YGcDdGUxbT6TcR9Fd/zZTycYlxngZVP8voXS0KNQ3UUtdOwK+3/UYw25Vi+iSqJJKix9gHQsDH2N
QsQ7c5mEpKkMxdD1W5hg3S8yrdtSD4TUmXWVEIzXvQtiwlwRzTwKJelym/fIJrtCnuXj14taCaB8
pqGS9E6WZvVTiXmQvFdmDunbpCe2qKKtVQFgiCbiVHFlT1qfDAb10CYiD8m+qGmUDC3mQhoD9Ce3
+nIsSGUxzU4WEYTrR1o7AYannJIOmegN/MWnY7mWm1Z4S1ivsiZ2hsTFxW+K3c6yXufvJJRZ+lRE
EclPb5exunQtXfNNQ3y7A9HJtyVfylwvxBMDmqWkV3+PNGCKADYgnBkLbACJvNtmBZdy+kHfZUem
LRrmvNn2aFdM+XQCWb5yASq99/19eHkgEkCqnVb2Nk2ESyLMLJVhfeS+162T11hq5KHVUqBNcVOJ
FtOwplRGjFsL+9O0HTzQ6a4uRo02GJBT/L4Y8hE5Lut79eUSn+SDibmUw2V74xeKIHs7t7XAtIOf
zB7+sLHhRZMXDhrzLnGOtJYJHMLp9rYt4q7je/U44N9p52hEl8EgTTCOdfzfM4wzb2YcLIApeecr
xSIbC3+RtIGNroe8vVdc4ELLPrjZuwm87ApcuXWCHOfUvmCFv0ydkmaaNFys9nJCF2ZZdtl9KCba
EKkpBmzejv1jL3LdyAgZLCsIXbK+gtHjuHrA/13HKSvEetYm8LLYTJD3hzBTx4wqx0TAxjtZzWyG
rovoNfvzdZPmWOzefj8UUbnbEqDb/ybEiaB/LqzxhBKOr2uXg8JDDkJ+AsAYHj80DJRPE5r5kgsU
SqcKxqe7Etf2o90TGC72t2/DfMIiI+M7u6fj4/mNFRko9aF9Nvu+/5iFQ3FptOpc0hhZV3AcOaLs
VgJlmCuTfnvwEOE0zsvsTdU6Yxrv4c5l73klzscFG98Pb3YFw4QOeYj4eq49Bx+TmXi8jniux78w
QUIpRyTPuUdYxopovGDfDsz137teXIugz2rRiupyCskrgpYKbsq26f1ArROqlKvUJ7v/6n+QFtxf
JRtSJL4RItAaAIKt6AuVGp2cuxvjAbTkcCnQVbVbB1uX58JmQxlg4qQjto0GHfiVAhaCQkOkrsN5
UqiYYzkb16Z3AN8rIa3Rv8ylIAHWZUyLRO9aMjDb4Yslmn2KTVmX7dLgQwt/JkVV1ntq0s58icS7
HXwQE5wQ2uqRvkCK+o4Zh3ExLvdVzqx3/4NrCBFsgHaskKsHonE7pALGBLBYcEpo1u0Q7nhjYyyy
E58Xq6NC28JNETqBDvH9VaZ3g4XeisSfITURJpx9pLxo8Frp7v7dMYiFz3h9VBR/RfM7aCVRDR6S
nsimtAZrfJXzOhF7Gf2SOaqWIo3yh80xLCwdWv+L/nHKf0MhxU6A0GqQNNex3emIl17PJCE/Ut17
xZohTaGvyTb4YodKx3PeyEjxMvb9KcvoqcN9STGcKGNTx/9XvNswdFaRTHHlrO30NLZKSyzNYNJq
3Mfv1LQLpadAji1gxNq2lDycmjgu2vHBrjHZkG2Weah71qLnABvIez6/vU6KyMqnh8vKWMU/rqMy
B867a6gb4+X0iN+5dBeD2qDWeFuIyo6mDZF4nTAKmbbHAjaBifOsozM5Ay3l1hJQeg4IamEp4uM9
hCi3O61yCS3q+kqMZ3bw88l44eS5497dDfkAOplia+sQ7gn76u5oyNzF/Eu+eTZkTai9mVPmgMYX
Th+gShIYEf1Ol+DmzTlKVTAn/qFXK0nm/iPbKYjIetBXY2X4VYff7laXHkl44yuSc2N4TXGVIuFU
IqqGv00XyZvUB2tW6YVnv0DIgYqhR7HUpRVLFRrfUTHX0ynWSp4uRYReZ938oFmPl/AHlvTRsyQT
KaSPyJ/i62TPG8xDx/3D/CIb6wgeJJB2VK8r3bzhmMEOKQQHwymC7gyA0qil/X4yt81T597oy7de
Kt9Jb44yJPVX5B4/jIHhyCxFstWRHfC1XURuvsyoDA/Gm9y8mdW8h9h9W5c0OrdAzUV6q/Yz6JTm
8q3a61I/iqtXijhiC/OduHF1Z6dUlCQdYXEP+bEsA41elG2lmf7JXpsHgCXFxyTMRXIKuALBh41K
waCHt+5+3JbQXZC13/os+wLV/BTeMAOEPaIK5VoZZ5bacx76zz7u3yhzvfqYF0pVl/bSPHLMMphU
CP4G0G3fIi28MQp3taMXxh0lFxrJm9QrSvNlfiRMIdYDEh22cMQ9rgo1v3sQGMv0igth6hUYH/7K
upDH6EzVh7ZsXv/CnjHDZVE00/A7WMmAB3lx5+WcfUo34Rpd1AFKX2jh9+ew1NLtesgsj8E3NPHr
Ee/13NgegCjOAN/dq8FfAXtFsoHnJ5xe9Ooz0TyigqzMC+D+Rntu2zufzHq6Kxu2R9J8k7n0noPx
UN5qRc73CYJ9XPHJ7VJh7g8B3YCBLD85W9rvkNLu8x3k6/HGGd8n/iDmfdFu7datFWZZnzXWwWpN
lc34WJe3b1f8pFi5jM10XApgOx6tQAhxyOYPA27dmrefDWs7obiUv+KXN57evwPuSJnDwBlfUN6U
SMR4ZrrQ7KSnxmL3berXySmkjC8KZOC77n2JUTaHka+gqkKVYqBYqEdWxK0FxS538HFlGhIPZj7l
em/3BI677rkPccdoFe11VmjsYJRFW6vW7Gf8NqLZI437elbd2Ku/3W4St9TsCkX1fYNWKpjgVQDJ
5LNUdZZLVAYwWjmsUrTa+IMkgArOHy94k2bcsDJgbPQtsyOAKJvO8VBFioDk2dGf2p144xuOHzCb
lfoSm/XASMP+39qTD6emE6MUGUla5wPRymNMUiI8x+50HZ7YCDf7bChBnx9JbM5GRC/Uijn4fnT+
vmBi0lheTtazN+iCitauleit9fR5GNDT+i7/kutMbjaARcT7ryQAL0Pc27YJ2fcaVXMtVDV9pyf2
NGQ3mBlvkaTYeF561pn7vxfgeCvdQlF72mDMSlkTMxqoaMlbpoun3GHzN/SGr6qmYHfTKtqsajES
FyyQPmnXiP4fw8X3vK6rVJpFEQOZinYoyveEOzdWRXQpv3NYoeT+r1D0ElB/U05g4qYOKS4F5oOo
02jPojvna3iBjMc8slmDFTjKAEq/uY9BC8jKRTnJ5e5S57UKRQxJK09XoG/lhE9C1yUGfOKYidfv
SePfZMdmZkD21KhnZa8eaSCxwDClmHi3cBMjR2HuqXQvAnd0lx94rIjKRHsrFjh0oJhmc7Rg/thl
3wN6/IAP9Xlc/NklKxlS6S4hfZIaC9BMWFX7WHpXZGa3tltI51k9l4qLZdP+RKHm7QOnDLhGbWJ/
N1b5eJLN8C0jpsb5OelD/FVKtfblbCDxQ/dL7P7G5DVUXzauNaB7kXy0skDQmEshBCDEucoUWbNt
zYYe0KLcl/Jkj6uSDWSdTdvrXlFzYi5MoPIyUdlS+dM+zuZIMNWu3Xk/fNl7RuDIP4n909cGWU0S
Eh8UDEd1nPYJQ0nBIWuAqqPcwGi/W/LZZgKSCIIO7qCIQrsoqMOnNJe3D2aQjYWozqY8cMCMFm1i
vDzs3p4aijrIJj3IeMwCtHBlTYxb76F9WzUm5V2OA6OrInZqGFdM2ycx12WdMICUcWfIPTqKgq14
Z9hlGvqpHCrTTZ8G+isPHx1hQYdO1ukTrz47o2teDXivnOwB2WQh1YKmvtLuNu1EAyNk9G0hv1+E
L0TI1b1QvuFqWnRtwGSLk6TL4nEsVRCTz8vOcIIGt1VVUutUjYT6WFlvwCb8LRIio/Qp+d78FiKU
4gAD6CqexHrTYidQEPaLaJW43+PmYmxa7vii66fQduswlcMEUt1iE2VciiaF+oe8q3utdHq4mdSc
YAE9/qvtxanCJ2NKdcV5dNp2avIecLEbuIHjS52E4BPlWaSV94a7CtpZ2Js5d0NTY/RSuyroqUTT
F2V/7qOCeid8EHW6p5Igc5nb2e8s64NV6CY0mkDjF2nC8CztJ1ueUu1hpEYJ4DYt/44pSbxTG3PW
TVkIQ7zWDxbj4j7ABGy86OpdkwILMGnIjC7SmS4jOsbQHpo4gflabF781AaA5wd+BAOl98wK/RQZ
Ms1tF7ihq8BQzzMsAKtPMFUPtDEMN+ChlaU7chIZIaSKRlnbt4nxHQjaFNrTmZRdlD7zfXjz/3tn
nd0CnVxMR4t4G/i5JxmUBZPvE7gemOLG0qFWrL9QwXq/LSOpYJdVQeIBas0J2ojve1/Ky/kFYntb
grf1q5TEyemsaN5n1da3AQnw8dOobvqbCT8KGCp1pp5jW2az/aSgPu84HCZRiJBc+VTo9DVopDaf
S7TLIwbPrVghYZXgHAxMJN1yyopjUWKhIsdCS0jrdGJaDj/wCU4OPyo9UfvoTIGkj7oWOcOdrodm
MxYEKTFk9+M8gHvwV43jLKAkOkZ281hq7yiINvnq5PdS2Tg7uZ63qZ1I3rKJN2h5PKMnHU75p5st
c4Qfr4iDK8ziAXi0rO2Nxa2PPmU0+KApZHlhxDVCR0406Kr7TRmZixNalRi4HvwLFF2POsqvUU0F
j3eNQaI+1GguxGDma4sLuvXtcADliO3DgX88oQzFaUQcZVovy8lYIJIoJma1UMN3iY6j/oofTR9d
bwHiu+wXboDOy3xIhhoBPSEDUfez5+O2IZWg+Q7Hhc/qvUp10hnldEfZawphHddKP4DwdxVZvGFB
0JH8I9gUVIpQD3bbcDuOGX0V9uS7KhJswoOr5W5wD0klj7yulFglTVT7FAM+0CE0TBC/vJXXFomE
6ASKo/VCZMsjPkhQKXWca1nASQf+In+J6KoPyOtSQ7BGdyzNZH1rcmRrGmmTyOWhW1YQxHnuXDil
+wgqj6ly3mCqN8ZXu+25c0u5d1gBqfx0IdWoVf0bNwk+vBIN/nEA6tNuPynjo+7SiEdKYk9gMuET
B0CeyffM2c+SSZVsm2a+d9C9bnzvEtfVnlJgr3s3rFgnhGrhhGQ33NQjQ4qg0jJQISf8ZJCQ/i+F
UFtlGvisi9oPLYAY49g0QTQQETxowEyR+bbPNbrT29ddVg8Xew1kp7qPbuoOXKiPPi1d4TIlIJhW
hRmc8pHjdWVVK753AUoshh6HP/SCbYWxdpBiQOzVaHSyizMjpoc/ku4c62UiUYQxaHC+3N4tmWQ0
rnFih8NDsG219jSfQtFPnwxROsPLIhi2bQAqtHMeWyxIIl4CkD0SI0c5xKyGsHu/jm+tfFtYH+mI
1H6xTyxgsLSipnVs+i0pYbgpVX7z+Jf/spVwtao2kiJRJjfVAQL7PSTOfjucGIEBYKFziz9i9dti
U+JeqNxCj0kQibdr7rhSdaS1+UBxkwfxRQ9M1ALA/N34ucfQCZHWXRYihHMnDp7X1eGe7Wkf1vza
kymZyCqfqukQYfQAGKnTSy24kg7i54YnNOSx2l2JvW/emLUu7+rhAB4KAMwWcfsGMDg4RcvPvcUv
VpG0gnM+PIkzNcHubQTTFx1i8mHzk3mSrhlmQsmzGIL/bdgOo0fHMFPqVJhAgK9UplyeGHvRqUdJ
4v7Kd2S4zErtLSho+1fCfsBX19wIHNMhTutT+Jbf8WX40oyiiTZXzgUZvU82jpQUOMBDe5WS6JaM
/Fh1hOb5Tu9idltX67rONnWxqrXZZDo4vxgKDsKNi3N2ciQaRPl4036Umv5qiFOaQO71OoudDija
sZ7gb5SgpWgX8lK0CVls3qQ7ws2Sysjzke7k20DkVR+Meq6p2VRvw8q1YQSkQ0pKkYwqOk5xTA6K
R6VMlOT7Awq4mvMh3X2JtZx5hkVX+8LPGwVAlDg7Ij23nx7AmRSQpoNCtKVpp58Y1BqBuIqUjFqc
n4A8YIpzhZHWCdiy+n/+1bwFFKtNmvboe0lhk3qdmt0fEjG4FZxstcytRX4EgL3SHjoRIh72EUdO
WCK46u6uO6DzU/Xn8uxlvsnLuBxqR7NNe4pPK7tDpKTPJwfRy6sURkuZqtVedfx22EDYzvyL0euS
pLKI54s/7Uu6V7XUgRguTqgWIOJ0vSyffUOGJbFsUfFU7xzzPGjFNVwl7aXz9Ww+F9AFR6mtjIS3
oQG9/tGQVwPWqp00aNmN5NJhEWSVmRLB0v+YJYR17yc69jikQ8cICxxvLayrk5u/wM5/5xee84ZE
Aq8Wg5RV2SEi8v8Cvrh5umw9RgWcgvdpAoNewIP21W8c5dX3AU+aX2oXBZx6+TOsbj5Ttu9d5lNp
dwQ39Xp6Uv5M/rK5BFYVhFiRmqXIRWNpVr6m2MumNuURKvuWl3O3Ge3OLiIEzwTLMP96ws8OxBOr
dagBlH+h43dq669o7Jms0yS+hUguZpoo0WF9lVmgfbj6ncM8D5/SGW7QTRtoP6nNbvCeP64HWu5w
1zI6PjAoas4gX+WHuwTNpEgKMqMGyx/KuVSqLm7cQpNs5IFzF3GXb5cWcIe1+7pX7hcCYSvzMRFH
WAylTCijqlfalCuGHEL6TZk4eOjI1/nVGALp6IpHQQrQnNZTM1Bcab5OEnr+53jTi4+WGzSNd2Zz
JBudRmVB/NpiUIgs0ZTVOR+IEKYBmFjyUGXcI+ddLYImvnpWwsqb8GeUl303PH5n9N3dPLXj2whz
DYs4hb22nrt/LazI+ynaxYnEI/Z5Fx9fCJOkE3xP74KlyYNt5mGpclhz3c9RCRIOF6gg2nVt6tfP
qgt1qmgE3tKB3gB34ooFQZ365YFH0AncH151vEwKnxEl4CB49xdiEVQCTaAGkjoXi5yrNFP8r4A1
RLIAG9XXwurqXda63dB/nBKpti5fYCezwo046jQE7uu/SH6vJlJwoHxTbbbbT1N5zD57EpS9wRPb
9KKXFuXaGdjDjYgHRfzy7djob9joCcg5PMY/mB4IH+owr06mlwtgBUmXROwY22pWXiORLkbUzuST
jbA0bhRHQChpjf1wUz7yeYKibNcmaxoqfxB6A/hNMZsqDF83PCVzq0iZQk6Q31YH/4qKauiM3sDi
rnJp6VqyWciaeC0El6GqbzFlQtCPhAJMeoZuvGUqngBL2YCywBu07IQbQS8CpyfnHrk6lhVSkFHZ
MgYG/x53nfTIShyiPRzYXH/hO60P29AQsioM1jNaYzipqNLU2MneMFBdgm6ErxNuZUAU52QvopB4
2Dm9q5WhowFuLkumhlOmk4Mk67x+0q08faTjTqZ+idB/QkPxeiCC6y1D+x43JcHeIqTG1q77NWct
VurYaFiTxUbUNRruUBwYVocOgpzA9rJCU6CF48/B40YdtPLmKk55d0geowYHzoHc0qbhJ+pwElqd
jaxsgXvvx9hPdZGmELZ/T/iPy4vP/iEAGalzDwx+9rryV/9dG3/XeUl/N9mIcB2H0qWwXj6bXrmq
un9DBoo5llKK5x0S/0qeJZIgjRsYDwJMh9eXA6MjRzVWnAvbvsugwdraNKwdaY3RRxws3oNXuKZa
XC3b5xFDlK9ryOZQMIxLAJ7FM67rWxSs0Wioo6hjd/R8I3hc4bIqJVKF0LCGc1g1yn0NF68NEQsT
8eqMfYS35IuAKSyW3VZROxdEPemhq+cFkKl8tspdUx3JUDThkh2m/rMNN71a+Q3SMNhtWzydmGAJ
TOyvyUS9ylZ4d33EpcMnfIvCWjJCudeM+MFHryKvEcvKuyujOIHvNAW/BHxBgxjIFwc/kK6nGziK
UFvP+frn2YSaRs/5EohBtIigIr7pTz0SLZIzy8hUQHjo2VU38xoIvYr8qYFmXpWRjh+QdlDUBuTy
1kR5ymL8NLyM8P6Jtb6f1V5vDw/ILpsqO4D6x8VTgN7iTKo/dCmXcqnHb6KpQV/qkaRe8N3DO5gj
LsAiw/EDykpjiJlDZzYW1qf9pyuh54M9hO86Z7Y+1HjX1/BkhrjWPEDWQekpu7UgMkzbR1IncEJm
jrGauDpKzUp1BG1Ub4RuBX3TdM/HkKSTAgmX5lQIfPaeMV9hTLBjMB2BW9iNtDvHCkafK6odUwC9
cQdeLTtHyBEDxPO8QFqtFH9r6HoaPHIr6hS9dQ/FvCzkGe2EC5CU78YZwLD3e2A6pcqIozi6ErWp
tS84hi32ey4cFFC45vJxkDzrbYeTqIztgKY6edDX8qNtY8KL/L4yoR67U7xfgb9WPlhXvXuinezx
2dBkaBW9ZO1HqlBObgLz+hyrfLmw/STWHge1k+tFNiOqhBoPdm5ttG9IrsHTqzr6q7gqh103vd6O
4Yt42QKkjnRyEjem0fjNlixWQK1WgcxDIOS0DWd8M5PQ3hep0HD8jVvUu9F3RZagqEWq9mhut2/e
mGA9SOPDOVoE7rJYvAz0SoNKGhSdDEK6qqsCFjkPGHCeBf0Sy25x3Q70r+P6Zjxlk40Nw2oequco
mahWBDFzMwHO5bXnxDwWk4bSLZ9i1hEa3f3n57RcgTWSz0tDNEvaTk6OSvyHRWrEOkt7qKYhnr82
Y++82v7d+ssptXNc/oMFh+ZdGjz6lFpBpQfK74b9D1GqsUn0FyKIEHOt5gjKHHm+qXAnAvs/2eYu
d0IYKOemTBf79VoeyyIwFoObPOKrmOrHtYmoGc4xnUE49iySIT8j8y+odDWu82js0T2J2SS61Wnw
1iUOFE0za+ABSQ4qHPrYrjNT/pyhkAdVe0ugen5Qok8HAXdwZEC4qujr5kLWgsa5ioJ45607o7wS
T9gz1g0+dJVTp+8K0S4x8+GiDI8B+41nJq5OYeRZ3EkXoPCH/oa7oqgjb5/4/C7SP9AOm4JZ5pBN
Kegae1yU+x8JyKRhRUk6OwbQorB6Z8s1jNi9mNvVXQ2ZBLhy2BHhaftoDuGp0FCmFy3DT0WTX1nl
2DFX88XL76DFuP0fmB8PmrY8Psam4t3uBpE7FbkjBNXVsqVmKZgebPNTxuS0Vy6DVYwXuPnbb9eJ
SRZclj0GuZtVv5oar9RMv/vb7IBYo2xydTlZnfzKzhzOuYqXCgUvUBRYXYKuz5b9gpknJ8wdigT5
7zi/IP06OJ46Ak4EYVrppVJewBKuDM1ZL29e1yKG+TlWbyr8+e63RgHo2geT1wm3M5Kvs8Xcmm6O
j3vb7/IsEDosDlBXsod9nTWzAPh7F0i9SlScNiyNrD6XQF5oSkQu14reNK2Ls9ru2X+mYM9vDoM7
6SDto+JngAs7r80lRQXYCPDG9ELShgBpr2BDLR/tU53RzA3fleuKzvIAeNnD8DawAntXm7WrU5xW
OJ49w9dk8rZ/2LVzeK10ahAWLP1+3P7ttZ5bSpXRYmgTrajsrL1SVnSx2xfLygRs1WOkWR0D8i2D
A+LBgbhAXh7JbvumHQ91H0fMs84RHlVSwRnwQAR2be+pPQpvb+IBumkUye8sepa8R6QVN5C47v45
diVr1CTOgB0daZ18/hpI/TSBWV1yku4sq1AjHqZdtPmL3bwor1xSX9Mk1RPDHx4GM6zXCTIcl7KQ
ZXjrxbk70a0E6/Jv3nh5f4uW0DjMYbjw1ezy6bCpPJ4GI68XgPu3FtyEBowf2f7nKumsd+xunn7J
4swBG+x0O9L2BvXPbZVgs27iSg4mUOahr3icFvCZ6Ax2PVfFpZX3ErIAVB2utdw4Fei6LYz96GvR
D9hu+XIDaBlcvUxf2o/0966sXpjOT+7Lc7ma4HC3RQkw5HGoRvcwrrYClctadtrYdYxZYFvo7Bw0
EZvivsRu+tZT7H0TBbgN899rnuqaYT/+GzPTikYxqKdbLBJOK4pTSs909fvndv9+q5/LnSqeKkiC
UswVVv1uFwQROQKOKOJnmJA75j56VFtIyjMC7mxdZh7v2nq/6B2r78+D2+rp3IRqwR20ch6xdhuX
4/u3q95gld7bfniodMQ5j2EeHHW5LzFTdQc0k30Tma/M8zNOy4a+bDDUqzgWdO8j98szuU9Ceb9K
AlpBSY10/TCokcjPrENyeIwJaFIO5eEGPABByUpZXHR+Cj8U308u3VID7MOtLROmeFgBCLqsLxll
LJPXda074RViBERTnrow4XTrLsAwJx5Ai4iNcdbUS6sK78BxRks9+5VK38VFggzSWCNOgTHJvUbv
6q04T0p6IserOZrg2wPIsMAQ2wYefyaRGFvi6b0GW8gQrBHbRWxcfn68Qc4zKwFLDaxMWFNnPIpV
FKAksn/tofiYaMJsGwXP7GFlKFhb3HTMiALmXC8NQ42naWkAXYD9lEoZzzw/2EA8brk5Wf9gAnXo
By3dlOMenIZR8e9NuGNS4lqAX3hU5y/iGF/IkmLL4oQnW1utyxaeNBs7T0OAsMp5A/MGzcRrwY5j
4LXcTrzfsBDVEjRxha2pr4Km5akWwPJuoFuqCMp0VTns429qC8O8g7q5Pp7K3Cr0yROhcBITaUCW
5fYRIlYFPnbDXLlrbRGdxzDpcxB+4x5JTIde/Yd15ud1NkTA+ShaPYHOAfJK7Y40r+QZpBwbB1rK
FSrJrShTbOrn1+oXFWJWjxGNL/H/MvAeOeFjdCTZo4vPb7gbFTzKUq+pwC2rArEaAhuf3BHbGxU/
IWmkzfZZg7aqNkBpFq9qM46w9MCqOM1fYGD1LcqvJ40WkK/u29VmSHKR+15TNgu9hHZo5WH6vJRm
HgczZibxgoOXjoRI4IuAjKVeqxkMtybGuclO1JFczoHf2HhHiwxXT3huwN4mxUau90DDYsIXZx6w
l58glp56lgifKP6L9FqMyxGcVCRqfArT2Q55H4LroA3ypa3KfDiAEbwRxcSXrP3+Tu3nkrzKavst
YabgGlUHzFoYr0ghyJNKAzOw08KCEeG9KLvb0MaS6grWxzLP+K6UIdqbD/MnyMKllwA759oF2y8q
8+zTJh36bnX4wDlvnxX7KqVw0anCcMWfQ9VFIosJyR2USpy5/V6wCr/hmW5X16PTb0oRa0084eMG
FlhbbcpUjTAW+T5u2ciHlS4St6Zqj9AklWmlUQpwor5UCa9Ix/tYhNNi6Fc8IXPfRe2kFDcGP4qb
dao+KPBDnU/rcxqx/n36MbHXqxJOwiO48lHNnnbmRW4DMvI57OqVgzToX4zA1CoOws3uVqkJk3FJ
qBxZUjWOxPWY0Ke9nrdVGo8rCs63EbPKeohTHmeq9K11F+swniV8tgkc7Fw6tQPTwvwSWndH7J28
hZtUUssJJjycAPD9QiKaHTATVVjggwgWvClXrO7WK3RsGuA1Bhor9pCMNz3cWTwboIGgfjiBOVYo
mRzVfy1mBM7IYlXeUwgVHlM70zuu8eQ8slCR/Os6mLj2ZHghVUyWBhD9JwvXGtzrAL1oVr/aE5Dy
tgSOxh/X8xVIbEfcYRAWLJKUKWMxx5YODqujytyx+uzQuVtfoP2vyVooj5xkla30m7RERQcw8Nol
2gBay9Xj4Fcg9Jcy+AXxDDaSN8XZAhN4wALMiKbfhCNHD/VszpbwpfXsyDx346JWSEig83Alu8rR
ct6BZNIWm5AJU8ydmtJWEirVBNAfJo0inw08thfdumm2CkKkzHeThh7G1qPQpxjcLcqKZ6KDoPt2
cJ7fYL8iz0xx17jPx+5Fttzjv4/gYG8MNJ6MmdhHJ0TAZZ0B/pv6GNVnaXWwR4UoL8f2KF0KAIwY
UgfmIymHcofPVgGxs4Y5pk3Qe25j16GExhOkkskuQK96Wsl9Xz6VFay6B/mLd0GJdCanXLnr4ISD
WDXHk/5eKJLCL1QHf1uwit9vlSDUtrYyQnqivVdyOi/GEu56tiZ/o14K2TQhUVdZ1pB2HN5YvhgH
ddyQvKdy7Ucc7Z3bcr47I7Dq2VW523eNg3C7gonS2UcBDK0FboAeKwJ3oo20PZjaZidx/I9UL7yO
uihh/LisZgno6uUgQzuGH2nm254FnsNFsecX2DbfVHHH4EtKeSK3stz/7cv1o4d8EgiIXO6H0AVb
R0O+NfsKsAdvqVTvn5wSUZ9Ai9Djo6Q5TQJrtIMLMJ44UtDpdAUfbz4iX5F6wCpVQJjmgmwYZWPH
OfqOZKK9epB6arZwYsR74+gM1FhuV/veCDEHgojvGoVkm8q0c6Wlls8h9sy5B1tohlpJAcHghXwI
6/2Fkte8pEnNyJDz2RjtqLKkDd86zlDeX5Q9bbJiNw58nARuHDzcYyhIrHW2xd3eKEZL8VuTvJM2
C1rryaWqZ3hpIQTVtHnPBwE88CwcqWnvE3Oe0zEBDZ83VfolatbHYJPobA2voDOSfLJuJJNBc60O
ltjnK0plh/LX34j7hWHn1HBPEpTAOJ9gBXk3h0S5gFnR9WCkYjNeQiaj44UeQ7FE+BngLLVylMUn
pSeoqmV1jUojpCTqb0HMFBILWR38JXVTvKyNBk9YCPsGtiiuBk8OVO839C5C7ihnBJ8+b/hC3zk+
XkhXnalEMn1Biu28aG2vuZOlmD9iTpFokOXT6qbeQon2X3jikrTxLoa9MUipD6hqUgLYbtMsPp7j
WTVXOpwJqzjrc9gEJ1hGYVs9HJ7uYLhap7E7HM7rFbwJR5jjqGMxYpxyPkK9dyOCW4qSBR+kJJg3
wL+/48/2LW7DzSg2pVVsGyFvbCz3F+lpNNJ4zbD2XhFG9LjXis1NIarW98hWn0bfNxbFMHRVofZD
fYAMaV+u3Yb8/P6UswePOesW83nP7RuefCjn6V5osR72+LvWwoeqBvEDIOz0MYFKvk6QjGG269gi
VdlYl0RvRDuNiCfi7GdKyml6D7u3Gbpftjs7MfJS0KqPT5YVyVQ7A728vBfvjI++T6ZCPlS0HeHo
6PlM6f2jlkaKecPi39rJiYtVesDqlzvT3cD4v+m9na83o8chJz44gsejTy9DimTy7wFNvpuQor+1
VcMovIpwL/ulPVupxVjRdcCuSeZxhd+i+CB2QralH5uSqZALqaqn5jkTGA+pLPV7XYq9y2dPmxve
9Ki7NaVgY8GNN6ZpSeIEJ2DJ2txtOnTPTNG47O8udSaZhMB3dRbfRaxKID/DwG9RlSmsje8AYLos
FxNw4GH5j76yTUvE8XKnrk+ipk8bAoeUZL6wH2eFeFcJsuitHjQibEhhSM97knPEoQ9n+EYnXBty
BiGGqFNw2Un8Y4z944DaIuGzrnl+kRQ2t7qWDvMH9mAp4J26DTiYhX6nMX7AnQqBwpW5cMmAxXeb
2fZ5MbNKzuCBRwuiw2xqpQ1LhvviQvCY94lw8DP8g25cQtM2TdnVQ1mAiLjQYNsmPz//No41NxLF
3XwiVtLRo00O7rPvBnhIYrjy62dP+sBRCTwdXNpnR4hPK4dFQwgmWsxDerqH/NqpuYekM/NkAs1e
3noO8TTis4TGkWNwh9en9aGNP4D1W4Xq+hzHeB7x4OfBEb0ABNrGcpBdp2n5qfV51OJXTINtIVY1
pGNcDzAzqnQnrc2wKwBBWYJKgSAYAGVkjRQ702rM+BDUHDRMc6NZmpKvp5oaiw8otZJljuUov5Qm
jPocktjgyaIFOlaqytohbgnvEydo0Yo2WsWjIr38KslW88ehdDKY/Yu2mi3RS0DXFZHSH+jnmmfK
4sBgeugkjd4NbyIpDp3DRbFvDttyWJn8Zj6RiYnZc8y/u6MvtQrKHUghON5ZNeTwg0fuNNYqQbM+
XTC/lsdWdmM/btbQ1WdvZzSbEKEQglsMwknTcLLnZ4KaL+8usIV0D+40Xr04qxgJYYlgj2kclFOc
DdOiZavUo0QkzE0LAQKiqZUMAjs7N7fPKo9XPCi67nE/wSqErettAMHBTpNq6aAE1iex+VRu1F1l
oBlest1LUCo5Ik5lwRI9IETHGCSMQB0C0YHMiog/qjmbJKRci2X+NW32eRN33P3Roa1DgwrtWPGD
7eqHBF9gdhcKWFxhAgrBF3z0Bw78rOnSe+8viqJFws9rJHqennboqXHZNEreEOs+rk+WE00QS4gk
9zWD59Xd8TZ/2p1wON2szLzExzjWA/o9t6LOChh8L4vLVd/ZaNNrCHIlW46vUpIpm9DUwRysOIZX
GxGwxBv8k0BCLkCZtykBEzY2Gh/4nRNuQywo8hyWN4aHbmw0Su4BKUyMwXEEKUcyYQc2xebL26zu
iwPpwEAk+s/Kl16+clYRnsTQlGaXtbpd6Ap4CLuM+5voTQs/uWlgVjeYyZOAz8SHJlsMg+vc3q1v
wmpFvz9fZ5I0TV/ziaDWAficLv2ApaXrI4KLuOW04lytbNx6GFTecL0+EtWRcCkL5iUu88lNQxc2
gB2jLV6Xgsv+M6d8/uVcNwpkmVEB5A4s24YmTNFFzh8u+Pzas8D9giEVfrDAidzvupZ8v/46ftiT
0pfvUPYq01RvxEgI7/Mq9Iaxvwe7uNw7xF6C9OYM9mfzTFV9o25wQKWikFC49f6DtXPwQuYhKPAc
N7zGs9MWl/OjYmC7AKcGLt24ubUOkp2NEgI5JUTgNQzMMQw0Y9O4EJ3GM8Uh5P0p2hi88fr4/yTF
QNSdY/TvoGCC+PMBMnmEQ/obXeoDXRDqeGjFj4y0eljGYxFdiUem/KgpPezmBvZ+lgbqA2HEUv2C
XygrVn9jTIMyzyeqWLzIZ4O+YAr22edAUPItIbcz/3IXpI1tvaFCzKCOJaH8Kp7MV8XnDQHlbLqW
pkW84ZIPjWyIp5IIkFnBEgr/FRNJjhlKckGO15EpUhYNsCVXWDMxSoW1Y3hQFUc4VUMOuSqqYPRa
g7win/dOeDf/2NJQQpmmhUVLI/1Vvwf3JuK/5V9LEu28V2PvJTeDk+pnaSaGPFjoGUIfMVTiTZQM
QVSP5yZo/bT01MQEiLDE+GieG8EYUswfh+CqayLRyYc63Q/7Yr/D5uU57seHENlB9XLdT/9jLm4I
ni7PsrZ/bGkTUPBpztFVypza0gS21nJctLY6v+rWuLs7OvQIAyHmwQdsIlCcrofahmMOFoA5HXUR
N2F3sdRoIgOobvlWyWT5tyTu9+QDskf7G0Gd5t8qkcycIue/Lc9lnTPRGpHNzsQohaxhs+yAZ6/C
z6Rcm8UezxPJ+eWoLuDQjnWRfaBX415HZBFWTWBYSHRz7aR8b2ZpOWJRuvv1Tfx4USWr4rbNkJLg
FjWp9VQO9IYEtvfjB30PTVOBJNu4Oi0AJQttfe5qqm0YI/vS+L8dFwjaYod/F57Wdk0rO8d+3RXl
0ZfFSt4KHyaAkRCzTk3f5KPR1wKrHQG0CxqCRH0bQw9Dz3HIbr1eOVhJEN2TJXjmLPVUmzi9yJtO
ZEYsBp/13bw+S/vy5jRR/ZLJBB3p/13S8J8gs7/0vbUaPRVo1TQzeH4ZlWPgoS6IP7JuzQVOq4h4
JZmfrRhTlQuOBIfS2b39FdhdTL2/4Zz+rW1YBzQEBKeLYtTZY3Z5n+QiDyCxzijcynEV5sws95KH
UhKbdUKZtd53OOGFvcBZbQzQpdbPxm2J6cRmn71Nm/t1upIuL+pSKRjVTXXqi/67C4TH2DtMF6JF
dnYvWYNN4ICnZ4Xvx7cQL7b5yfOHXfqzbFY7JXggEQr+oChhHF4xkt8edTYWFo25DIrO//kEJHux
UgqOwQlBsHOwKuObhT2jZSDD9n2u9C7kLOgsnveyye/GA20t9CbO3AjQtqWFv6680xXx503pi6K5
y51oQtlmnSeIwTNxBFzS8PCGvS8w37h8i0Q0a2k9i1QP1aiHgQKrojSQCtJ4Gn2qX8t50ZP7J6pi
+iruvX7bqPs8vsHaBfczcJHaB/AXMRKF0yS4YiKyIEXpq+s6m/Dnf/IwsID+jWcCtVRqvV5Iogga
TiLA2x8KJTvnD6xLyGTX6gHfgxBUZk0TWSPHQi28ukDkn1BwSybIZ6zN/yaTLt/74qQ/ajYLPJPR
67X4QXyzEMoeNmwKN/zfn3cCAW5Cvf+7gYUtB6+pzAQObfmOXLrq5flhPOZFng3v2WL+VyzQbOnv
bw6GQymoyyr5kGDbdikrMcC05qcKCpoQ8T4yvb/+Bdgu7LBVnp/OOU9xXx6veCDcTzBwcT+Aozxk
WGujlvSxiw5qiR3dzSq9oSMTwEoiMvlv+Wkq45LvtrS1+YLFdeipriUtZqotneFmpCFndAs0M6oI
a4KAehOvWV7TMQu5HiA1ZAka0myQejwhuXi4suk4ZlaQUuZy1p18YAt6V4E0Bp2srH4TDqfrDRp7
Fyo0eM5FL+0a55Br0+oL50ArMJfc01NpuEI9avtCWgk2iX0S4gkCfK5100ElpbSjhdiRwReH051N
ZJhZCFmDuK2BAfCKqK4PrA2wHgimqXHv0npC3VTgNvDKz8rv+4X51IM4549H8/6AhMHLWO9hpMZW
0fJxPznBuRhgOoUf7LrTwAgLfDRI+NaSsRkeIDq9c8Z8pqD1QGieTavPNNljDW0JNDfGcqdZtEWj
tst07xF/nLMYRFRY2fCXyq72uWZ6+U6kEdZbQt4XrlNTGgB0eai1TdAA2z5dSpHlPagXKZv0eY4J
YSCaZVmeIyCy/oviNBoVo+pZgpiQh+1ddRrDZBuScS0/c2y7DBkOsKk7bVfafSBU3s8K79xNcbQs
yc1YbgERQvAD/sooKZCLBJTcSLVMdbvrmGvM2lQT1ZqSfZXxfJFC+5s/D5+/wR6DkTnWX9HNuI2W
jpZPiRj6V8CchnBXdvb5QniwAfznL97UuCnqIxHnEwaz2a7yDE6H7muvUA8qkLVjqgWfWJ7Y7mAA
8gJfA0TM8FOxy3x0PB4OADjyKTFz9l8jQkI8uESdCAoHvana4Kcoyw1daGHLCrCNzDGBWQKtKys9
Vcayd2PMqsgGriGqOcNX54vklEwsa8SCzTKRUJT+v/DkfBiRfQhrbhJWjwkpdCVi8SVcvGxWgczU
YzP4VQSBaOkJ/ywQqZShUNiBuXxwDgUQamLN1IVeWi3tNaT8/aUvhG3lb0LvqmeHEXgDLeeay+YJ
ZHuxri8uwjfMIlHPufm6sBuEaPbBPuVUG4EJlrDQOlkP/yj0yBP8xXAdFOQY0NiXBZHwkcLhKxWR
HVr3O4pSbl/p7kwnQfoLOrU2ZfpCi+9WKwK9rHPEDCL4Xn06uaDRQmF6SnIbpEI8zJVMBjN74zuC
/StEfR4eVItv0+fH7sKEz2pRdrrfw2xWF41Jlysj0u8CuhKMQ9zSKcw+1eST43lznHqF7wLM0sVg
K6j1OuHPdDzcotoRG3l7ZsLKb8FVAryiwY5271Jo43xeuvybADZRtPRYlmOjicU4yOa8yy70hkrA
bgMZK65GU4CFS9FTsxBv99R/2xUQr4cN7iboyt2Twl1lqr/2GjT0SHD8YUaOP33XDqnNw9K3XzyY
vR31IcR5Pk5/gD1nDgRRl5eaYzcbNkwBndsDs+vZTtSt7g0Hs3eH21TKLDMKDsh+NfFOoljys6MN
/Qm60az0cZIV1NbriUEm6eK04pot5ynkujahUtDA19DCUxaI9Qk/FWI/QB99jHTyRCNv+cAogjD/
203WiTDos11D9aFOTYmNBc5COnN2LKZon2qZKjvRgo9//mELsQok24+isBAKPpR/II+Zc6U8Hx7N
JrY4cLo1AVsQEOpCb1+VyHm7eOPh4g7A33w5kWYPPtQOmYXLuMXbH9Pd80BE/XADXbZQNy4B8Qv/
UjzCzy1NzIrvi+HRmuYBZzjvhZjSccdBWC/TSvcJ9fWhniXssacM3zl8XGkKhk/e21HqDDohX+Nr
RiIwtetxSuaN8IAC1dlNUlVpoIRdK3LHrPPXMCoGX9weKwH5eRDBsGBicKroTtv9mJa+q83KNY9p
hAleGVTJ9nbS69zxnlLguvpYOp31NkcsQm6o3ee7vWZ884Yazshl3tBxxj2l52h1MWdwBoPbrU/G
JYFrBGQWYXgOlJPCqoOChWUayYSseVbWdVKGbdukLPYeuv032gRWVV1vXm1bjRHvbYbQflvj7TgE
VsddW1CJ9XDWwfMcWTxr2kPE+GF3d8kEavblCz3L8HQCxDp9bgM9DiOsa4MlrC8OxG9xhf0InT7U
9UdKB2kQqsMGv+mx5P8hl9Rht8xm/AW2Y493MzMbePWm8YFIcrDDg84ib9BaU88cR1LaVRg2jpSR
fVAUnAnFFWpN+/hS7+rAHOSdDKT1aMHatbrZ5uUGejHR2uyBXSteehynxRhSmo9jCqu7QNvDBU6I
QvLdSBG0wD9DE9XF1gN+HoJHR4qdItdEmbkqRygCmA4UAY7g5KpRcXsNfqML97eU0y4Blap5+hyw
njQVd/zoP7dvmQ4M8G15BQQzpfi41MavPuIUMsiUjbkz1CZQwVR1Dae2Ji3lUH+4jiQ2QurXoNZS
cDYWU+q7SPtx7Akvytb8ok3dWYqEqLZNuTrdGka32NlfEbcwqtQRc8VUyPnDiLcwgEfkGVXLXK+7
qB5+JwMWEwsUefALYk47Ng5ZvX33IKIQR04IWlGGqPM4LdMjUKIo65/8uBUbJU52r1Qf4comuKHT
dQPo2htiqHSg2TYQVl/8NTG9BIQS41scpWCxwanwPrPbhFzjdJvvlOWU47VJ/hpDGOvECST1UCfc
t4p4ie2OCQEVBtZwQPBfCtVRmz09phI8nb8tsFhwP0vdBebF+44n/BiAaGmkB0SP11kW/Y0kmgjC
3dEY+rCF5zjK832ln4CxUSg/Jo8V31U5ZqC+c/T87f9YiaLCq9NJjEflAEdFae3DhW7tKC1mlvPQ
XpB77wbzGvZiQRllTNPx0BtSTkl30z3Ews49HcrFNTa3XuvBqYJD/QuPBdsQIIeEC4+ID4wkytFh
8Zzs1NXWfUaCvEibqlr+aozxjbzYb3KNigWDTLS5z2PeO3l2rqwhXeqJUYcDeOuLPrNQqWiTFIuv
2z9S1EVGYt/zndrX3g7hSSSO0xj166lv39UgluVAH+Refwm+gQPCs/B01raC3xso/UHZ64SkoUbb
TdBVr3nKBTOQC1VPLkDbv3oYK4WWR9bXmd67+05s97T88tQ4YNxgqpKfDUgRWdaimVp5t9eq53zI
QGNf4LJ4fRHyOPN1gO220iKMw/o+jKKhDR4Pinb55IlwnAx1JOT7vkGRJ+Rq8xQgcq7AqWCcZ+CB
T/2bAhAF7WF7uw2hwLGbbriMqXaD2YlEnwIgUGrpcoHBHCWhfhKKxXno6igHHrltLIfChP8pBFib
6vyD6gflJfIXcVnfhhrF5LCXeLTpTzt3TUalxL3F0U66Sjuf3jPM+yCx8+72UYuDvMMrhzg1KVYj
fjj4BWZbBMG0TySpQpaE91G3wSdM2wdIREwi1oQCjfFcrdbYI3QhsS0LzFvKQLIuYrmA+xMns1dT
hVCKvzsWT+/L7lJ/l/C3ll0dXZFa57JV9/uBTUwHO/ZLcaeh4wfLb/h8mryBu4SATKBog+DFKEZ2
g6LriH7S0O/KUTfDy29Xs05ZgwhDiuS2zPj66Z7Tto98in9N+LHJZRQCfUspfWbamJYMorKPDrnI
BKNrb24fL0+x67WwFAshzu6Xddt2tBuPf/zPrBIbxmCv3+bKH48HHCOZ3wIhAG4AWaMn1Ap9sYfb
3i8m8GdAw7/m1Y4CzrXO0pvNzmE0qAG5o16abDYbjRR0rO1xmybmANVPrU+pHipJmFar0Xnn9zP4
eBXrFr2MucSmxnEwwCa+HQzdzSSGcO3UMcOwQBhvxldtT1r1TQcsqXraJPFmjH3e6ZsNz05xIaHJ
z6dkSuYijRhdZobb0Pxc6onQQ9oM746qM/JwuVwguazrqi5dkp64jaRxBsOlOyvDysEmHVEoeQDi
XQptnuqSeACk8UJbu9qMswl12gq/42Nlrfb3u612rpkTC69CW9FF8vWDCwPthJ1838FD7kSS029k
uKnU0qrZQ4+kqbCyADfpfbOgX3W2ta1SOiRGXLlKfi6HGS2D1i779mYM3O8swLdZp3JAsoaSrKZK
q5k0C0aVx5qrrWo6iZT/Tk0D1GDauJ04070e9eMrN8y9c42+IRAQB+F1tpX4ejLoNLxwJM5Yu8st
4ADTxy+NqOfk4hHxQhvwml83O7GG+PDPkCCqQkTZkeSt745Wa/nvSdDl2ahnq05PUfpScwvya0IM
L4e8hrxU5FgLXYlLSw5wZ5V5fwgIgNRSkcMa3KRNKz4kOkvFZNW+XTVFE54TbOOskR1CsVaOIerW
PbVUQ6vRhHrjyJUo51iRQpdEGmc3kjFUb1tCxcoD4uNuBq8BW+T5otqAvOwTD1qlZgzbUmFfDoRk
0MXCcRddtp0mOd6JWwOzxyx7tm9U5kcvA1QRFdBsQ72gTLrtbjZ7T+xCwWc9moezbbDy6kWA1kk/
gvItE5foUCdSEPRBePk2IiP/pR4FYVddt8RixpDdValVQf1+CCk4gKWapSxtNOchkr3ubPzIUBey
pL9ddk+CrotAx4T23IvA5LJIVaGmWfWq2odDtQHTiIqRYP6aM3wQQLWGSn+Y1HM2aDrHFpn4hynG
tB5NGbLgY2P+uot7Z0NEjHf1Oxr97n5g2OUwoJw0sebZyVq4lTrLRY5ZHvGRHDmX/QEnLDBII6IA
0Lx4zxAoS7uIDzmqsNlmUFNz4lO0zwcfdr9XiDzSJMXT4i/5nV2alh/6n9T6aE4I+XD7oUQeBl9Q
gRjlofYRw2nZseX8Rc9abqLASCm9rWKoccoGginndSlS4Mkmnbqpqnd3Zc8C++Afc4Blw4MLQnCC
hQ0X+NS74xSX1/vVWAMPrJE97gv3D8t1jKEpArlt2lls8K+HzCa0IzKnJsvK++32zu1UkloUtJ3h
8x2L7Rw84pbONkhlah+DzV6Jw5r3M6yrfYUc8vguxff5Is+8qGpxn9JIrzmLnPpOQHdGtwolmZ/K
XOezzNPIACm3xvmUKJoklXBWQS/BDzrU9dLoEWg/zVHr5zzs+Qv6qPGNOZvJ9D6r4FN9d+OVAVXg
An2G4FRXL47fOng0bZ93ujCM4A8fRONN8UUJ+7iQWSaDbOROxmBFY7o0a2CqBcp/ARxKwEQj8CwV
zBAzUfwxIERJW/8F9pPEy24JWuRE73WRRzxi4n009Ieu3iXluEJpetXTUSz2N5j0CxOysgTg1G88
WuB9VO+WVO90niFN84qAGRTTePv7Oyw4Fb1GF0PdqaygxMQJZPCHEJsLzMeVMUtVEFMSPEBceY+7
iezDtad7QW9/Z3UZCpWxCpTrJaTZT05EqyODTgrbIJzrigEYLJBuumDOX+oUZ8mQMS8QT1vxtdiY
1s9SS+DxBByVoPRmxllkY6FF9ltQY5chz23g0vBUNTMmLL0koLj+3EYQ7zfdq7CX0WKjJBeoBqLv
rXoiuUGFMYk4fXXHBJ00cSL5ZwkjFp/KJ4Y5WyXKkJQUlsTx3UoBxEm8LjVIOuYjY2iJ+Ky9N/In
LpxWdgziOH4HdY9/Ev/7t+K5k1covofUUudpNxGHinHV/uHd+mLRM2xUL83jHKLW90s0fDGxm+uG
pVWfDm0469DKgGdsE1DUYOF5bv9S1292auR3hLsJCRLzp6CPCgPySKPUiSD2HZ5m+n6afK05ptwi
75apUHxK85pN9Fejszcs+mNtZpmTWvhF7qZHCTe3lB4EJNZ/0CHwatDNiK9yviKwiYr4lyrd1+wo
iXpxs+Qg3HgukIwkNbz6MYYdn7gk3TKUkEjjnALAQJER3g0l4W1Xe5p/0lAk37Zr17opUjRW8MF1
AQ9I5SDmOOH0s3efNzAcDwtodJjAP6SAdX1Z8wh+vQh42PZeeIGlgwEX9HkSmB6K/UF6x5Jaq0my
DbewA1A5PP+mTl0aUAHxajChg9bUereF4yDSksBXzz5GkuNO6zr2QLw8xWtJ0ejK6aZEJczyDo6/
tijbguumUnc/RQCy4k1cxapG3ji55N62S84visqk4vapVvCwaJafIr4cuCiIaJiBlWOSaTDMj8u2
yQVcmAqgA8h5a0nnxYAnGVLA376hBPScTrVMtmzkEnyI1hbO25Lg0YFwipEBrCwWdiXC10o/tvnB
tYJAMlV8G8w151K6BvhnP4Rj8cxkBd1jlvgGjUHFq/B8iU77cRwqICum2nqjLWIoS0Tyl43ZdN3c
s0fx5AVgIkypo3Zyb/AgYjU4BJUwfmKqK/x/rgySryTkSz3XmUFKrfdCePpeWmRsSZwXY3rHDcFw
/0XOzHlq+fZqWb/CkH9vQQy32KAfeKRiQUmF33wK0tC+Sc51T7MwCag3phmYzG8r/CD2JueXev5e
2zKdYEnS3nXs/ljHoq5OIvYhBKGCveNAYUggev3E5GP00Blp16CJpn/3uwxoeaPCvLHjdFHln143
U6w/aGo9J4jgE+i/59+83Bjxcw+FT2ajUglhxFzADwMlCxS13EyBSGZ+RL+nMXi0lCs3yJvGxWZV
rRQhNb7pjRtMJavOfciWV++YqObqinOoeKJahB5Y4JKI/kIsEkeFbZ3MWVVSDqMw7CvxrRLs/68S
nkbfpEAV12zy32onQTajea4jWpECJzXFCLy2W3EANW/it6wDNOVMUtr8H04geN3fO5Eo2vLcfrax
wJDOicF+5ShOGp8py4tdgQ6OZO/lL8Agfg64+gnBmWKVkXigc4wmMQEiIuDo/Maze51zOnc2QPYU
OU5DWQ6I3yeTKYgIDMsS4fr2HIsxOne9wwrRUXnEH7HJgrug1LGOxe5erymQfxv6ZNhg+CAg2zOr
kt6pY1Ey+VwOFSLibuMQSHvpne+47euaR/fOu+GAq2vl/GltrEw7WZlGLjdD7E8MCxxqNW/razAc
10GMqqk5+zEXt8d02ScFqomNXr2e7jtFPfMSRz2NGM1sk/sncRGR1mKiGRS/q+JM9Vbrw0Rif8yw
ibk3z6y7NNjhia2BCBpC/uzZ9oOMc8LVf9y3W1dkR2kcMIIxV1ltN8EdSYZvex+d3wJp4pkHAume
Iiv+r82hmHHW8xOwq5iYXtteCK6hBxqgxvk5aPR/XfCiq6/HwSBzLwuL5SZRbCOs0hzWfLBWOf7z
hGpq6xmVQYnq6BMxhv1JfPl/Pq9yqSixkxf1JFcmNjdOANG2t9TzbTeKot9p/y9R+ON/OlSU6t57
W92aXNmsUG7d7hiwT90HI+3xigg9Q1wEehzXZ7N5+mpXNSLykZE3eh7rZydf9NjCoV72EdNLsAsY
T8d2NxLpAyaactBL8pIVxAnEs1i0GqXoCD81ZuXvxF43k85puwUv9AwCGOGVVSqW6xhve4hzn8eW
ALPDn+nUrH0+381dHZGcJvB6uVUkuLEUU+LpPqiT4WRIvOH+oPq2QV4i88xOINyodJUGIjo+XJqe
dIB+raHDaaSgNWhn6MIrdiHfWuDJft5cDwqFAMzhJ/6P4CWwL08EQ8wsAg1E/LZDOGewLwgg4Hhl
VhibtG/ATjolZBkBg+h0MJMzL+3u+TqXAK4ZvwWxOJhTwMFJTNN1HhbYv5HMtMrNIx/1yLvSZFgz
1HDsnciMLqy9806IHeHuf7QQK1ZZdxEqEieEJPhfUi51tFYIh+UGDk17AQHvZv6fZwus0YFR4qoX
mu8j8TXklmnG2H4e/dgTnjCIxESQrCQYwOFFrySQ58AUsj3m8b211wsqx9SHAK/XQFrYETiiwvm4
Zb+EsonKpvio0PBofezpCcJRmKx9HJQVvQ64OvDLb8xq43444LzsEd50ruzHHTJZGZvMUvwalmQU
YQBARy8MwaKSQgBGULoWnSqb7HyxuwypRLV8sU7Yi5I0JZGwdjMrMRou662LwQUOEJFH0IPv5sOh
PxDzNO0OpDqkmVb8pviKqxY6AKWk3L2wwDcv0X2hA3Y5DV6wEj2dPxTeD0NGPjujtoWpCOqjKXlR
TjoONPgoyLyr1d4xNnlgzu6JMljmkbdMlyD1dlDf70ybTvn4Rh56PiUnsHrZMCnTziVhlqtq/pjB
apsfZgaay0U6nDubXNP2z1a+p3lnR9XCWXeYshIdZfCDc/NN0/3x5if8Opd3qLG2/VZCSZ7Y6mWW
K7MJaDK9GCUuElkJ+7ABTiPn9lEwf5SoTVx6EYgqBllz1dwxO8QOXx3sMM0dyFnhN7zrg20M9kvq
Sq/SBEsyLvTf5oJTE/SxPSfoE6aFRaYCkY/TTC9aBeQ5OIM1exu2C5NwjJPEPuED7LbZ+HCD6l05
mGMzvYePC+uAhQf75tMRILXWnXBLGLUiOfekfJi1cvsrfL1E1D3SidrxANngtuvR0Jw/kicYzloP
mFd6TxgQ+o6AuChXSPzgZVlq0zkjnUxoNVIfOtJZXiGGwSHLZHCGxpCZQt9/Q2l5ZmWblWwatf6a
cjUCyq3yMAtBhPT3t6h1o/+2KulOJ2CPyF0wFn8G3Lx2BBzBnk6ChShA0VDblqFlcFcNukrlX1fr
bn2Dr0x7mJVIcdi6UQqSVqOlk/n9W7dl3xInzeV+N5aHEOb2v/A0ycc9w3DfDFBl+LaFlOUsNeST
4GMkdZbkOmCMBQtyze5BhdppoYTbQC/r/FpNJmmTUZqxAkmJTzBrp0E3xuRD/a0H3RAsU110VIoG
yOf6q6lhVEHte5IVEV6bvnoOJq6k8KEhmSaxi0U9UTR/rWKZgMcY4stEP4/ikIfPkBETUnt9t5z6
EzlGkHeuQhEffnumfhQ2oubDrintf0TCexnUEpJaO5WOhVisuvnmLI4GKOTAba86ORzaNS2RbYor
MMwj38wADj0HDmTnHdQ1K61S6/h9Oy7pExtACDxc0LH0nJOPaU+Z/pq+G0OBr/WlC7V5K+oZYEA3
3nRhohTtHgmvYVmkeNX2AfnXnh2M7V+nsyCIbHnNL7v6J3N1dishG7QGE94VphPY+Y1yqLwO6zXw
z/5xwJzGvVJI1woWbjODYnjYIdBRn46KqYaG6cjKiMxHe99n7D/scx51rLD8uEGxgt+Sq2Nfe8hA
pZo7eg8BDmiWfn9QQ53dyZ1J9vNAM8DAKGJqlUEytNecKocpCGNx/AJ6StJDPedBcHEOWIBOMom9
AZp7Rdndm6vQ6xmFth+g8tQAHXtpXkjeopPN4ezgTJcxsB+DJJNtaFn8IhJTJADKI4HIUKYdTezr
IbJJsqzFjwF1UCJjPrY0QiU3cWll6iq0O4rgvw9Lv3mCsCPSvxqBwFAIhJqA1k96QnuRlvj87Hkk
Odr7m+qMQ44sxXErpSspC/8k6t1kHwebyUN1/YLx/SCCOFldmCjsSmx7TtaRV9DdKuFycw/Sx+yH
MHk7uBBNtOVAlhJc6XJWqjdxDaEYklwg0tZXeVD+n9pY5P+49akSiSxhqsj2oOsBF4/LT90VeD2V
j1bmSY6QY6J49/P5l+UBXQ052uhf7RCwTwTqZakebGKQvrp3B0GwqgYQfWFfYDAg6J567uKtCJTS
pTHUytYu7sBQnsxrFYfEBalJ2v/+oHIhBR1okSitFeB/1YjGMaGkhGaAGfa7secM/ctzo3LUdIZV
k+ggjgS/IcQ9lfYY5RQDE4Z6AfUyhFtbKINjM20dTYXDyUe09KqWX6w5tEo5xe4ClXnlQALjM72A
sJBPJ93l+kP+vmEDk3WQEkAI0HLtCPrBQiAV4KoVpyYAUm49bwYvPKh/dzKXOsKqjwRrd+WyxnHF
Wn6pc7hgnHRPVzGHDds4b3FGZB1CxZ1cPRg7UDKZJkNiZpt5QvBEFMzqRiPOduMAvgkRCM0OUbvu
820eX0ysAHl0V/k42vmyhbfrLoEPxMYu2uiWGLNVtTrfpM7ROdaoBuayzJW2oDGKnnYKibGeEwR1
1dBwVO97XR5/G50L0KYbhzqHZ8eitrGt2xrfsEGgI9wWLZnYLXcS6B1iD8ixtCA8Luw0DblGkojx
LTv8CkO1bRh3nVYJe9Vyh92sI/kgd6XAGLBU630j9X+5Tddkc5Z2wkN55ET7W9G1H4XCoiUBXypw
SBAd5xpAZwYdUta7e03P9m7N5CzX3hwMS15FvOHNCuDAtqfffDaNGMRPuu4MNIkXb/3/0DuLmolZ
/oTIiqguzkHPk+cAEixnFLRdsjuS0zglVizKO41n5jTmdQ6gq90p0WxM4MnWlWR1DcJOsZ889pi8
Ax7Z06I9OVo0Jg3atND1q61N5LSvkj19XqzUrfCDrX2b5x3Y9Ec37EMHCSPZxzYzsWVaNtoWpXxI
+U2vTJe7DSGODDrCM0SRCWf7uFChwumZmZ5nHgnBhWu3yFklQGBpQe8MDSVyaKIj8o4PNvz5CBVw
fqE18xvVKBUqK0jUefuroodg6BndKfHi07K++awtTeU1a5ecQSSunwKoECg0btwMqdsz8+Lq/mrw
iwJZavvam99e9oads6/zoSiwHPEt/tV0e+9RbA2j/7mXWz/uNyvvPJIlipD/EJlZ9uxlz4yus09n
ECarqMTUavM8jAZha+VGMVm+cMoAMVRIWCz5+LrYzKDQ1lNlRX15FWoB66M/PuVtsJy0iPtcMvux
TTOPPAXzOLmCbhxRDPkXzME0TV0OJb0fQGkUYSToINTsHNk775vVPQ6bF40J5l318INkas+e4GTO
uySCaXO0bT84aN951Y3UM53G6yQBi07xDtLTanGFPY/vQ41kWrfMXyTydRKTonoziHGfRoEP5ywH
6SMzyd/b5y9WXfWmvC2z6OtkpDRiXzsdTf6zKtlyrKJmw8czZ12R8MxLXYzn6f3IX7bnwb5srXRF
boCU8N7tptb+Imp7B6WnoEsyytcpgkWF9oC1UHjK8f7DSNgznN3dvHiUJqZSav0TImbyMKANc8t5
8+CHNF9wLV2NX/CaWzV273I0Tv7qRglXHCY6QtOyvlY8utjlpz1d+ONcVdWQTu8M72COiZ8glvYn
k8uMoODIZCSpBhH7KJDu91T1RqRC06hVayM0wEAjY8vFRFptT682PU76T6xFpq84pnW6AxpTVVcN
DLusoZ/Q2HGcPrUUvriF7NI5Jf6ozOmyWcaE/dnh1+z0wKUApWwxlwr9XL6p+5fKkncynoXFmB5J
l57R+tHj5An0/hx6mkMfVC+Cwis/UMPjrLdvyHrZC/H22oo1eyz2kJaBe7sCVa/GclhW+hxqogzR
GSSSyQlJcAzeg8rjhIJGnP+KOXYNAmWdyXVmR6FeDAO5ooMJI7l/8v/k1OZ0TFBvRFBylafHVOmu
SVC6xJt2+3pmcnXHOT5YLLZIn9pdqLsaZX1+m1RvMO5g58OBYhRJj0Rpsw62stES0+MdQMgZxXQX
2LQ/aPBOWEjXgHLOyK6JH3/crCRxug/AZHWgFowrWtutNm2kFrpQE1ef3tY+0L4lCCVlUbMJVCNd
Ue8Rnvr97IJem1syOTxzFqoo06jemQDYssYzeTj9YNjQS//N6bfqAcUdVlzzIyNA305kutQxmmb9
yKM5Hhz3GHx9U4YyqwTEi9D8XyceOeJ0TIVC0jKnT2ysyvXrYV2FYzCKfUaAyUh1c5UnlQWTIfRW
QURgu+Zy3PY7i2uBqb5RFm4dxd7R8qgVpmocBU6GoMpex8utji7n4OQTEFzGlF2Ylca7a2WKU+EV
KtzdOHdb+jMPIpfVX41xuW1MmX30o91YhVIlQv7MDly+dNVp0QLQ69qaLWXp6rwwt3OinC03OTEa
dLEvXjoljd4hzagotFmRPWwqlnzHtTLBUONuTN/hdRJzF9Ar5pM02TWpjN7493BKd8QAeI7iNgAy
V4DwyWXXG42BLHwOlCKfvTtPDfo7IaG8v4EXlLSDVy6G6XRaXCv2Z+RMupLzZ/0uBFPnvdR8UFDn
zSj6rkd861Sou5n37lMHPUPkBy9VJGt60Cww8A16l79HnfnFWr/sP8QbaHxwIhTb0KpLdA/JLdmt
aZWG67E7eHJmr/Mkujy7l5F4PV+GgChI4Kew0ZaU5P6OyQczaQBHA5q5Z3aqtKe3HmUd+oeTAWQ+
OKCwYhP44fl+XjLWlFzMbr3aZYGkbncryZWaFm7wUkjRm8HgbCjB3cyWKB9kQItpDLWWdvL23y5v
8lpaBmcWjckNbUbF9Nhd/yYSmf04fcxcOX83Uozu72I4ZF0rxGjtwxFOzmD5ri/aFfec9s3fqmrm
C6IZGxoj+hdoGbn68ippn3t3m4An5Wb+TPJtfTWsUSEVTK2vIKLymZfehz7ZxS2wrHIb7ACH1DRC
1H3VMwRzUM29VUGTXo9mThE44sshYJvuvzePc0pXKeSvcl05Ng+l9ueMjaRf2PhOdFOq94xxXhNP
2FhQgv829SeithWhNjvCLdF2qalC6RkD9vy59lT6uDqOm8O1V/Cec/J0EWsTUtkYTQByzbsm2t0i
mKoLTuNpzU5vzDDbikVJQ/Y4v25YCh+YOHmpK7Mhnqml9Mql/BlGTV+2h5VWAGFs4ZUh6R0DOIk6
4Ej2VrDGMljU81JAmFtbUSPgB7eW5AeYgWbXVSKWEx/4XYZLu0fCjx75Pdh5o1hIaCucF4BtDeSd
PElMSGUc/iWVptKhDfNSuxHoss7hQGg1yQCLCpypKFjIWvngRxlkjJV4xGZPHf91XTQPqrF1Kn+R
K+kYQc1Spw==
`protect end_protected
