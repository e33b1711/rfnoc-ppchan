`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iEjoYdpoxcGKWZRsp4oxv+EZEzUSeeVTTkaAPRciDJnSfbEPLLKYk8WjFSfy5JIAkkCfE3q0nnVh
qprJuZXAhg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e9ONTVGwRJLTG237UzoAJdABQ5rkM6DnHXF/sF1/uVdMNCBT3fG0w+FoDhz8kXvk6j1iqmQ1uNA9
MK3DBbhknUW2va8MH0azAZdGR6GBdKzGZYE8QuUtH6j5P9PkRg4SZTnRUtqO2jJ8RZLOqd+teMAJ
E6o8SRMPuN9nafQBGnI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S88fbr3xQzQUmg9JRSN/GAfY/ZzDfycX8xGttAB4ljVrK+/Ud2wPf2T8zdM9B+9tK6YnyyKTucss
I0M7aYVXOoOJ619pvkbCvMkvYup1ThvrvX2r1cAwS+XWnXhhm1JU8GTYUnkF4TqjhaH76Yh5u/EJ
DkQ8dkPQEL8szNDBY37WanHciweZteIA2EQ4bs3Ao8G1B1hOKp3n6vnSZxJXhpdHcqkaCUufdqaM
FrinxwWhd2b8vF7Oemr3OSlqM845sfCrMN7jxAAgHLAM0MSMgfKTq4o8CRsTHWQQzAOPoqsx4fzF
mp1LX8/oirmCsufy9CIJjtJkQ5LMad2v2GOxng==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C3UZmTnXNO2JOGNm/uXG4U8HlhAkjOphRlJCOT90GxGNHlPsgnu+YFgyMxXFTOuWMzkcEiU3Hua2
KsBVrQZL/9/nADC8Bse8IldxE8W/BOHRy1TparHAlHZ8f7botWVRTz8IoKsY6ckC7flbSTrOvlyz
+5nXc2aXR+lsQkX6n60=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sRP5Gn9NwCjZeAz8hSSnN0il59CdKNjwYzXW+sllZnVXN/N5yMoHSeI89GYIqBSGSsb21UVo80nC
dBxojivyuUfqpZS+t8++R4eRbffR31bBUrrSVg5OosCxPxSCHv5hLr7xlyVNtUmQRka6Y8Wnyy28
blH9if9JaVp2t7EInlr0a+t8wf9k5dP5A+bQyuu5Kp4nDwYAhs959ckVmufTJxVslYSH8VAMtrma
FNvPsmO3pTxY7bZ/PEIDLrFc0xA0mvB2Un0+Z8TOrxywRFfV7kMy4JyJOJ3WcAqeFWr4la5LuoH9
T2OLtZeG7TTN6g/8bQwzuQY2sSWtxugM04q/Jw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CTYJN3IGTSMmDt4BcedvsCRhsSnxHT0LScK1/qkByuKrhygZj+r7nAppYsaK2eQJyT5AZNIKYyYD
PwobzSlRvdtK+Ju2XN41o4Gj3J73RzyJgni8RHg9cUcf6lZfEDC0NJesqtbaVfEUy+LRJkpkmdWU
GLgqGSDsnf7fw8RjZ+9nxPuUCJgbOp6zwafzrF4VL7aYffqyx/M7Z8fxyq17ga7TU/prOzR35ZIk
uh3XOxTHUbGjUroCj3VA6LZo2TTNBh3OQZBRdL6lGNwRqc3B+I2bfUE4RotHIOs8kqNPu5I0o5CB
G6PFbQ/NHr/rSrdVyogIDq+TPL62jsSQ/f/twA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6000)
`protect data_block
+W3fXb7xlQiLxlTFROgPopkt67KDN7EWIVMJdJIfzuo0XaPffin6eg5gOandX0bh3walwFbFMV5D
ShzBHn3bQqn20i/sR8t0zuJ3OjLLeyROq9BMZXHR42G21JtR9G5+9BpZ4UI/5q3eVI15aEohhktX
FnA8yiYXKLoPsCwrOrbiseh6gXCgMY4YDxSAmryCDffWXzb+FlDEmpanv1fnRV2U3YaSMMx2sM9E
cM3aG9urCt8QJC7MIkSbDqL2NR7cX3Yr+CpTvUsGlQBPQWZgF1m1zzcz3CI+4R4COELQ1FJb6vH+
RIJhENByRzWY7PoObBRpz65oicGrob9efG44et1R5fctVySAAAkMe4VA3PgdORT3bt/MWxA7l0/t
1ABgTQ5RXybS/7TvV3LcBPDX7JuSQHYXM4c/7Bywp2Pwxm/3Z5GszNSlKaBOXnYfxJ1xr7117/Rm
tm3l8Fu7yohansD0b8BzNBJ+B0lBQ/ejPEH8gWTHVgZK55K7WTK6SzJuyjs5svxtlt/M5KD+nb10
eveEuThl9tMVVVZ2DRsy8PZJ8BuvyY1RGFxJX7zvOV49miRhzis8/P3vKs5RBfunVCpi3MGRl+fF
HTJs1Vfq3TTCGF8MODhYAHwqPnswVuN9v/eyCd7RA/3OqD/lghY6zo1QMlrA9dpFcRf+gijcjOTt
opAQPldE88h0vnxYvslRoT10nBHuT+Uep0y7+dDgH3k2J2OTz/F3SowuPGq+atX29xjhwOr9qNXl
7+YJ0zqp6yHbyNZhpUZCTDoss8UlT5Flr9Kkso5ilNH1C8YxDqD6HqUdS0eCYF8BaH80Z+bnCqli
Y9p3a5WV1zw6Vx5wi17u7hwwmpiNk0BGS8VWIJ/mTOOlZilLwAtiXfC+ZBiPWOA4/T/wVyL5x9/8
IivtdByOi4N72sUS+7dZWNX4ifVxaMTaKmR4BbaKBlRTmCQvIN4qsBDK6gvnvVNh1sUIMJKQMo8n
CtRjY//ho2I8pzVyv+nJom1Vb87t4wuACo0NXVT4OF2Uy2PGXiFJcnrVUYt8UmBIJHQ5AtfX4q8O
TjgbU+l0VKqlljDbRiAFM8s3Gn5N2WPJ+v5g7sGaZnZvsolF+8Kc9Y6RklahIaKUkvK4SA4LYs/S
S58zOrJMzB2JwkOWoH7RHffPsSBWfkVx+br2xzCC6J3IQ9ouMvtSqRlQHiD2IxuVbwBMHBIboGwt
Q0jao9ZJ48i4cziRqc4n31WQ1MmlCzrkoF6D+Y2xqgmgwy2QXFa6SQgyQgk2Greipsk1jxV1zVed
uFdy4w4CjSBRdjJI1C90+7plQZ1foWUxHlAMBO8naRC6rhh0CLyD5ej/zDwsyx84id0/IbWoUO8y
+CdZq1ltcU5Q+1N6ywfugulQ0nXkv7gaDCKmlaWwL0WRx7OjK6ION2Xls7nRDRmQhsL/jMlQxQkd
7he5isYJsB6hEFsEKVuo3UXz/VpAUG7b7fg2TLHFwHcz4TrQyv4yuzPpbl45frhQo5KsMZ+X/GII
lwF+5czFEpE0y8QW0aGcTVrTwxMv0NHvq4NmSIUyKf+USb6yUYEZQIh/jtZxo0zdUqHvE60Hf82/
VeJDFLDW9LNmfVVQYXU+nGYhsdQtOw10cDrAxwJzX/ItOXKSB2p4O7ir4esxvdngte8VSp8GAfUC
GdHlBqyrM8sK3YaB6rT68TRB6NhzHuT1WnCYa9HpgrAKVcbizv4EGqNavmmiB62jOnIE+5Cn91w/
R2E9yDZ/qInbzCDDeSkqjPgQGG26mVkVWXJGYqCKGdaMMw45k+lH29cDoNrr2lefgssqgnAdHTmJ
WRH9vEipN7h+8ZqgRjrVAq+OoKSWTNlAoG4m/gZ8QoH8FeoRjhUi4UejVNo7MzJEWLKsWcmtvEQn
oQYEAv7cib7RXTvS8rtFRxyxjbSYGPw0041TnICrR41nC/DjoDladxYUQ4MBSnCXnTIxl6f94ZPh
THeiUWtUVO7Q1sB5qFd2QRL1+EtAsrjdRmsvYii0j2x3wtYmDrGVtoKFOI0JomF9iFzkYXZ29yKq
eIJYNLB3TP4HBTStE3AzM5YbzAolCr6runwvNXZCQA5AUfvuVVwjYkFxtB//ltbiNsURU0T7+4Zt
yQHsy3HFvqLfQMrLfM2WKVAGzDJ43WucHZ3hzHCshVwkHsCjbsLwnS6YYUfmbq0WLyP/94B5Wb9x
bcNUSJZ5V6tUvAexnzNufxsOR+wsgClvFWHrn3VdkTs+XGbL3hz+skaKdNzv6IMDkSkdNp24o8IV
W5pLJO8tpz3R3WHtxB2bUy5wxFR2nRfkSqkOH1Hy4UNS1bzn1JtbJUmvdorMXZHYSJfMIxX4AAfG
EkX2sZRAThiDjRP45CL2yfQ60P3iKFC+E1DwXYbibL+hjFLD0S8ldThCQS1LxvDhimS8jz2UBOmE
7rYFLU+o6n39Ap0kUh+l7Ly2cDkNq6eulVReeJurgiGUszzMWz69w0i1qx/LhK/M0TvCFxolpOmr
7Nzez8KNinjSQQCmFnJLqBId6ss/2yYGh48gnOAO7Tps5gAC2FhItRSyFo7IGqoLTdusMaQiiSCE
YFS4AQ5MUQ72/AUsJNY7U43XQj9CWufmKYV0s2U98pyH8Sp6oiYbEgxnopXvW5+RyimbX0Y1wPjU
bVVOdKXi2+yII3NjMVfMfQDCtGRlDg7RcPIEfaqtnib9VJdJzestPo471symzqdEkXcUMgGT4kAY
TZgBjz5Dtu5hfL3nIt0yfCUYW/BXYSlmpPBVPV3zWwrFnAVq8B9uIh+5n1BXoWeqagX7um0F/jsx
1Uq3/8iDrWsROvwnfpl4hghXr1A2nfrdvd1op0Jg7YBHSP5eTpR/b47SL1VILqyuJ4fKiW1WXV+D
7Ss/Av9Dwtocts6AU+km0k+eoNkBz1Ix/6nLLjmqbpkZrJzY87h+RBf43E5UM/1b3FmVo7epDxYu
V78vEWcYY9Jj8eqhDyGiSASusiLItlqCj3eu+d6/un7Tm9gbGKCdSQjU6MVSSWwvJ7SiRELhW8Ba
7HmNyKtzH+lf57BG+IaRBs70obEtRiUyyZWGo86lEAgLTpJMfy49dUG38vTBOMEe4ex6UXUpkVL4
+WW0S04bBY5nkjWVciVQ8t7um9wHx2YlZ9eHXhpW9xWQtCJUAyi3uIHD1OdQ06eIL9WJs38RVtrc
PZu9F3cI6WJVh8FrKx8/YlweNI5nYXbQ1N/OBV8b9EdbzFbwzHsoo9JbqvgH2tAFO8TCSUQ+gT6R
Yu37pcPICPnhnoXmjJDFJoUwXauqtfrXDJRAcnFqNPJZ1KTyF5b4nDwaw/kawy8Wxfl4Gqi+CIsJ
JGGoldlm86mLrGCQZsZ0JrH2Dce1O0zh5RM1bhjLIJgcVCbmSDDyQClmjxdGTBvVmJ2iXzs7/04z
nd7QjYGXvlu5z2WClSeQaRIrBamNWQYUKDdnIhVBsbLFJWEr9NlRoqEaaPQW9d3fLzYMM3ykK35v
1gXoG158RCDU15GKFspkSYaFBO+05FT2Oddg7P7lMlVvVzIngquFO/cOgFbKMs1IN7jKkgU4MPsE
5qCKisyh2P3BfLRjqLjSGZkcpx/TmlpBoR4XDGrxDweVlZpxjme9Ffk8OfMoorZbXjGsO0CK3C3R
VQBH0AAno9zyu+u8zflb/QNdjYlr5u+lcKN+CDdBW3HSs5NEWHyD4NBa6LOd703edbAhz8Ftjhrr
701R7qQSOk1ySDSygmuaN9DJ5z8V2E0zcRUBw82npkLFw6H5S2nuw5sL16iqygeshZ0K477sGSNo
/yr++kHBYFkIxgQKh3yjzPL1QP8GmqYWTPX4FfBB1JUBgtt0FERNcrT74QDzsYCLr5b1Kq9Ii1JV
+hHAjnAw9ap1xjTs8+BN/ihX9m6JMHL1Y2BOFkpEci7d69KtE6ZbUm2bE0UsuEfP2o1nmAF6IHw6
fskBvr0UTOOSN5CmbgXYyu+cCDFZSGVm2hmBOEYCmSESO13jMMb1XR6tzMhLBfY+5uQxffnWRdF2
6roMgsgXOmo9pAKMY3DY8cSlQC019oI40igaM1hmXQGMFt+An4bQVBedCuUHHinpbzKcUO/eyMl8
nyz3N17qQPWYnmqE/ZxoPXmvrh7otW6BYHkoSxjN2u4JtFuaYy5vPuEatnEidJ/ZESvea5//Bg+j
AFOKu5SdcNpJznusUmMeW5km63w8pS9NMqxjfuX7VZK0IaihNIRyX+hkSaKkLdP4/04ZwdqlZITL
LR1HBY0w3UP2frwcDsKMhl6LVNY8lCU08BFc67ahB07UYhZTD/AbHGCVWL5jDlrnDfTsSmS3jFZ+
osRcmo3p5pjJykEYlMqi6bRN25XeUzOF3AbVpKTB5xD6lCp7wE6YOIjwTW3MJW0+O91bdiJG0DhZ
UxHcwnHuOOpUBA7vumA0/dFHEr3TQGsHNrMfiz18rNhkOsIykKYiTcPAXW41kw3+jshBBNFuLjqo
aN0I+NBQQNEQf5MJZ12qrDaUjF2SaYQj1wiBNrdR1epsKByC3EpxuLztCF4P3LT/cpVLlljrvaMO
AjMyLG51u/eWh3AQPa0QkkozyFMudW2OEtg/bQhFaok7IpUImeF4z5NflcfGYv2i2GhRohd6/k/H
DB5ip5pnreSAlQTkYTv1QM9hXtap9TpiaGaEU2cCUyKYTNx3rAK+hYdP5JZ64I9mxnZRKrlUiTN1
FfkWFZAQP8nK8283V1i4AHLzf/cRK514t4ndIBOXBB59xkhqCpfzzXv+HXMWYeVVphAx5ZVXMWdx
lWfl6cI0Q3r/oP5YO2VkpOSoTnhTzJptCuPqPsVDK/QT2ZF2l6MaS6H9tc5zLVjdNWA1UdO+p3O9
8Vhifp5QxDlH5xUN3fPF+H5nSUvgSPKKbKscMsXwlHIWNythE2GxNzUwwfHDUwDS0gvldzeYS3QJ
1kjB/Uhy6s5xQfXIxrWOQdgbYpYDKzY5G8p4cVddpESL/HSgE+M7HlofHt4uf7HPeIRQmP4k2eyf
yzAaGJVP6w5e2jFQCBRnn96CcA2aMV7BKdOZL+9OTNKo/MY9/RY6xLkdfedCP6IzmXlRbK4kC453
TywwxGntOQbCIC942Ed80jy0qvuNejRa1I/hEsn878599j4qBGyExXxdk033SRoNQteeHbcjSDHQ
ukMcw4mmAqxqtNnqmF/D7EvfgtQM5Yfukl/r/ioBUH5b3LJ0fUwb230jjc9x66Namvi4rXONs6Re
jc1xVq93F20WBt8JXtQWjGz5mEyQNE1qQ7qlmc9e6mLaziDVn4BqevehM+q6KgDv0Yt6nrFv55fF
JiEV7dhFJhBFkpUYiOu1ZEBSRQU8hEvSg1k5RZaBVzhVfUVvtzjOmhocc4rtV9DWYE1biVgOuYbk
3FN9EoTq8Qx6BOgYzX8b/plxOBeTM+f47ZAFIovOrJARPPPjMp2bwE+bCfBQKeLNskhgNmB/KheW
QL35nX6UcxBqmcJ1NDpaSZqXXsjM0oAp57ozr2nWGSiVZ02K/1iUEbs5d9w3PYRXFHgU/BOFMWe3
GURutL+eXWOO9vZQZwz7KRShLCpjPjM8c8IYEdxWy/GowAo65FzwVgsUUC3/pJwaxxwdU6q0XILH
FKMaRJ20A7NY3Rh14Hfgo6LoIVLYScny2aRALvypqKsuXOg94It/J5uHTtbu4SWfH7JRXMIHs+jX
ti1aOJeADdM/rl9OiBhLJv/zb8V38EWsLfULSKEGgbWMh4h8x4QVUZAidnrnuDJlwl6QVFUZgFjO
VxVMasdwWKQboAjDcpY31BAhMJIJw2Y84MRlCS7mjakE/weYMA8Rnpvob24+caGnYtjRnZusF7MO
2bl0rVQHe1m3p3mJCyapu9C+wzUNwDAQQKSJRnq+udrqdJ22MKwRMfF5x9VHHuI7SYoafvvOlynY
blagg/aU3oRzgF6+gBsIEVGgSKWDXBVVlz1yoAl1FSVAfTuA4d+tkeRXWk35ZEFd4v6FTXoJ33kt
mBWIi2ud38x/FsFIeEd1JReYY/jHlHVyp0T85C39WbF6TXY3TjQLGIj5krkSm53HsXxsBZ+cVhuz
PFsEpLHr5YtokKiruPFOD8trncYITZ1mizARfter4hgU0PPnxsQMX3QDqrpmpQAkXhM/zAKQFLkK
cbMbkFjA6LyXVc6He899NJFkTAAyYYdQjIh26iR9UQyOF81KEuKzuyeA87QRVetgFyg4hOyGHSUO
QNUl5f+bZnZt8A0c38tGu34pSHyiedJ/gavQ1fQHFQ/rV1wpEcJN5L5TkFPuPVaVXpkEd08Yq9kB
fgow35jBO4xPElZV1EeWEi05xvjqJWOXE4Pv9wN/+eWp3V+t0Lhjbi5+WXcbA7KVKQ7hZP/UUoEJ
0r8eKU0cGfbOWj7nf6wZKIg4ODkaG1wt5VqGtYVSj8ZWfGj+bzBTXB8aOb8CvDQuTmO1mIMR4hTw
U1yTTUIOWl/+WNLJba5Zdvga8QkrWH6IUDYwDDBH6WF5a18DlJlLZD6Nkz91pxSW+U8uqoDE+1hO
V37g2BDDsQGJteIGvP7hVgvrACHEy/TonRWqhlifMV6NxuWPudt5gTcvwVjodGO68T5a0681kDtL
Un+v8Lbkmhg05nkd8m8XmBeigq8x/Hq6GLYXZGxm6Mvj77qXVemS7MsfsVhTfPTDR6qulx4TJoBj
/GkDje0bFv1jgn167/x00i+ZQbrBLwPFUu/BnXdaiEcB0KvBYvJo1BDzhB5MqVEuxBT7wxyPqSn7
gGbUHvewgPmXXt98rOLycvzcpF+WDeJV1uxKabMEEoRYNNzDbKXEfHGyqsvjEPR0zFGegEyzUSin
vLnmreufuU7gE0FnqnsDfHs2cVzsB30/aJH/55xO6QdUBcTbXdQC2Acbfgo7Rib+VtHfsbmokOPJ
iz0pKBFYjQ9Yowp9A5N9mv2+uO2XTOI+IkKkz/amKWpstzrw4yFN+UNjURBeRJOa3ZcOgRJNHlZu
HR0O6SaNuPj8Gk3sRUv37h4b9MVyK8p+jy8bEomG6PNBHrvEm7zk55YBjNHD8xNx9zRPs7u+prmm
4YAaD8/4QW4HhHFk5/JtA3aJ7tOZ0rUxGVriOL43pjxIO22iJqwsZRiZAid8RV0Ibi3mrH7rMp4Q
q7hfOdVgGQPwp/Jis54e4kfXe6k6SLhhMV3MVIfXclDnpcRkNQXmY8QHGQYIulek9yCv4BELpbGN
wDnE+VPovdfNdXFoDeciCk0uAxf6HXHFt+5t/eTx613ap3A3+DYW9oOgE95BDrYzppPd2m1TQjBv
fz/nYopsP1G+4bmjTgIWKV4TMKEr4qc78RAdK72frUuLM/4hJlz1Kl4xJxb9R3SOr9zLJYsUCQid
58VJuUGe+qyvb3YLjXohxNovjNAeyGuKROQqtmNwklJUQyOWjZvaKSC18JqEMgGc20jiTCdsGoLM
Geb3Iye6a5UnH4P8/jpPl4QKq2pBLjJln+MdhlGl4gpdYnLJrV3cafC06hP3FpwmUhlHGtio6/+R
Uhn+6YLKEEymZX4rfnhuBM80uFkBrErn/N2xOaD4S+hTVdaPhf24cloEid3p5oFXr5WZbP+MIfLs
1qe3FXIBaBmsSls60SdDjv2wbVp3zJijAvrvcPgbvrq19nfPgss1/Fd/lCD1RLl29ar9dsy+c+w7
P2YHJwpp51PIElT1chs8S3EAMyUs6UL3Iqt36lvMU3fDHJy7/Ndb9kyYCnHVDWkxpi6t2OBfnQ54
krxChO5AzeceT99Dh4V6q+9XX+rrKW/ib2kj2C5x1LoNlus/Ods+tCtXyk6203Mt+kXJCY7XY2ja
CDSIz8fKA0OXBiEuvE94gkc7wBSIiC0nQ05lKHGu//aja5GW6U9/HEjcvhhlGGDarGX285fd+VkA
mJerPog+Yo5g0oSipfjd7RA5PHOeqCCcEMNyOLql8EuxYpt/854dnMUAmvmAhT4ANuTx9r5bo0sr
JsUkWJC5zBDcZLy7ZSoV
`protect end_protected
