`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Z7wtcnqzGEl1YB6x0obJMp/QqasJsGXn7Ovi+vN+pcuf0Kq9/fsmmFzgWzo2PqsjSidw1UDyOfwD
NJMcBJ25zw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TvSSJnXRDTx95zdF03mcP0Nw12huSfiWyui0LS6ZLFjdeo0Pfhv+n2rJavkC3Rp/ZreaLA0XtnLY
rJhjf6642Dq2FQbT7plurVPc8cCLm4aS4orvOJ+Nzv3aRw8UF5gqSlpLdnFsbBl88Xgpjd6DN6vO
hB6bDI3GujhM1pCgEuA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i9/MXTmWw68UYy7En5jmBz+lfIjUO4OkqvGPJqVxTaE0GIBqKseUmxjxrPZEAVLfZYuLDjtGTFFV
xI8JQcBkrlZaCzf4bp78wrAh7st2VujUi9c4ytSmo5PmsSz2IO3gyOw/lOqaYo2YFpHI3pC1Yzce
4JwoJCk/ZVSUfhO+DVAi3y6r6GvPuHNZspcnpolDnbiRZeUrv9gaizfK5afE8qnqMWS4DaEb1WWO
UUn5hZov4ELjgOMCXCjQdEpsX3C8e01yvjD1mK4VZU2cYi+NmZqxOQQy/eDOu3HY0/5uDHqtLGwD
WtJ4DbYcGblTLikRa+3ucLiJhAbNKS+xw/0TVQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zQb7Yu1jeLbG2rH/QGVJyx9WsuufurwlisJ4N5lJs19vc3mFW/MrorYiDBMz8/ZeNbWD9TmO1N15
a6qUT6qawxKXFY/O7hZKIjsVohny35oYjiJp4algKGmiXY6c1zt3ZUbi1z2OccTHSFNMCGIVq3dN
LkJc7cXJl4LqmQqm8fM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BWFO4UcSG4iRfIccMCi7CSeEXuKFkyVMa9CEeM4t23gWAKDtC8AthCnilNOWseLqMDNOu6AchXv7
NevbxD6l6gEL+jczD0lFztdQ61sDcwyKJJhwVlpkP52gErtKxPBejGg8ab9sUv0wCsNt/uTWexST
QKsCcBqIVIDVHJ0Co0jzjBRe++MWa+LU2y94SbJSv5sVC6V2FsumS7IEwUsBkZAbSoMVtQLqsxsy
wjYp/6QVGrRwn0Z9ogpH292TkKG2w9+RUC94IBRwaKWouN4C02nAXuplG6Y6ARvX9ZdgeYTIcXfD
jD/V3wYBt9PMFHEorbEmIj8ZhE53TeoSYVI7zw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gEOGo1TNktG0WMV70jAzFa1dLrb9izaZuDIzmneayRNzUfoCoWD4OzyomeOWT5R7QSFPZG4Noz4J
Kdkl/VhK5dCyS3Hc9BADzqjmkJBLWiXlzv8f+s6Kz4tgjnduDJ+/lPLhAT8YMyAg8dyf9ZObsylp
JNrUQmdVoxA9erwgasXpvfcCnUtC9SGhkD1EYMQTKJfGBIFWcdu6HmtwVZeMry5J1qFHaNKpFxHS
5on14/dcR+rD12bA8M39SnAVl/UDGnlxm3861bAN2lblrWDD87a4Sh1OHsaKaQfXcvLyb1iz4sgC
sGooooUTWU7Lk87EQwMbun8Mu6QRxVWR99hH1Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 93184)
`protect data_block
n2C2vFxAn2YB3grmWtGYzhlTf49Tc5ooKSNsPtS0wTcO7fvPx19gFv8+Np49q+7StcpFwo8yhzvR
0DE5/zoH4q//vuT2BT42WOW97XgN4KDeIMs64axVbhEm9OQYXtkCIPu6JF6PK154Z/Bggg3MYcV0
+VV6g257dHB96+GwKWHOIN00mQ2KkI+ozXiE8u3C+An27NLr0IiveQIDaR7PQcCVFNmmmvBV74R/
PwJiJc8G0QjUz603wLa0ClQ9g+qqyyu4fz4EWxTxNMe0dgnHaYXPEqzUL+fBg8U4wVbmThyeRgwS
Q6afvt5KlUvA91gk/S8qz5Rc6lVUtvZi23583a0FgG4TvLcvfs0sdNByFDxArJNB27fl6wBaolCX
/QNEZDGn/EIXhF/q5WhXoKTx7Ks0ooWY5ya6tUqusIhMc1AWjXD/rRed+xmt3XfW9n6MryJ0wNEe
9Th0OghW4az32aJ+Ned2FjFXHIhO14v+td2gS1fUrX6jwW8DzBUu+rmk5V4aLhJlDHs9jvr2vy/o
2996noIHf5bZ1IPRCGPVFF5rMgDGVgjoTaRK/xJXEN09MxpzW/yLuRfil39Y6mTfZ1DmXMuKhYMm
mFkZr7wNVzDSlwBtFOR7Ig13iq+bhlhXEnj7IgE5JIShTeQ6KYbyTonBTloXmjJ+X4eDdXI7XVak
Gn8dkOP2eRQEF4UjnkF/o0gz5ue/rKJcQtO1BREESY4ybuebkWzt+mW11hWvbSnMcoeXy4qsvMMY
duDciCk+1TcqxiDqC0YXKF6B9faE2xw6A1vOHMpzBXue/phzZ5rMjFe4FhDDUw1QusuBFMxVFjAv
bMb6gkBLfPwxSR97iQEBVl1f0OwPbZBp6ZQL6DfCm1Q1T39JtAwT23qR6bCeTLz+/oAzdS2EZn39
sGwg2ACO7+B0uzwSATqSpyx/+hp+ALdCEDKevq2cfomTwJOH6wEAE5zHlAw4u8TRUSt8BfCYrhf7
Lfh64prqLiYUjaBBhVwm4ZUI6pEJr38VHx3PUOREOdyzWl2ikH7ZLqbZ5EaEmVLnSd0i+qWFfJdy
8S1IndU5QnOIPWwyMwMbocIJiMIHhKzYb7dmHJIMuSRcyN9DPHcv9Wyoxt87b/g6GmdXUibGLIVD
CrXvTdpFzYKV5Blz6oSmJAnaHS3ZXc+GKgmuqvRNmf6h1VYIIqqbDYL6ayiuSciLGF8+7mBj25/O
o7LhcE4z14DxqpN+haCjoJ9PmjaMUGVMOSvTfOqD3qWprmglUmBC/f+LgO1GjsWUpqno9R+BgBAj
iRs4gBC3OrI/7hoyjy9ih5ZjXtrv3zE8ASnCM7xx7YZdl5QMF95O8LycOsf81n6p0kOVg6vZMZl1
Pr17YSwLGho+v0G6FAovDLHi7OxufOlLEwEC/DvNPX3FFZ+bd988/t1FqGouezhAno1rWkoh6zVD
VN7KLuKumKtaUV+uzXvAVYgX69yPBQ3OYZ3qoxQo32K2QtvKML1wzzSmyd269hsg3ZHEXziBu6Me
fnUBshRDV6ApE76gv6Bn2FE6AhgQSkCKcYgLahNTEWMPuWUxwc5Et2B6omKCRv2XkaVQ9/CMea8Y
pzMU+qz7ivsK3k9h79+UF8/qqpHRnM8R9tgM8B0gmWPnetCvDCd7yQh/tgFvT9741utNszC8mRgL
LO6wzhaNuSossf9MEqj4bxH2Hsnw7cWcnq7ubcSLiwvbe2peWbgo2TbtJkoa/YbzTfzFSi2zvqAG
9Ei5TgdfYLOOlJbprW3R1XNOClLF5CmTJyQFf07t2XDThbA/3xaZwX7BgHkrNqlCkqLLPjKACfM7
L1yqYdK6eaT/72Xlx/cxwMIGGH5GOsj9FX1m1iuUR5IrI+oJghm5Ld8bqJ3pC7Y0ydIV3abJzbIJ
57IWaB1MBe8+9v+rUlRktMmv2SoQZINZkQIwKJgNspmZO8CW82C68ncVpXcfEOk0DyA3GFTjbxWJ
jX+Oge4RcwQn/a0N7RCoh32yOD8JwAQGwScM2r0vJVkGMRgkEKY8k7/eq1BsHCXspHAkCccwkg4l
+l5nOLH9cbXwuQgKVCkLOFdykhBrgFUk0VrdWmsX1aAOShsi16ths43tSIoXXPNi35l+qMVKx2ps
njKecMwzinIIq1HGrqOQzeloBxkCeyJaBTZq4Gevs3qo0lzFfpxEaUBgQVIzeZaroEXfY7SJ2NsC
UhLbIxZwRJRGuEixHGSSQjRs10zaAZSBahb4duP4neiDzbzKJs6lJr9Bi5eT9szV6UZzZkz9qVwc
F+z58BLa/2MBFvpSlUvUvycEKeVgyiKJQ3fEsZWeYXVLJ6GgN9WTNooGNovnnJ5HWG1HaLeZgCqH
6VeUthVnFYbCJRiPV5sRqzoNc07oGr3hCczF8c0QeZ24aLGtpsEzBVeVLO+H0IODGKsMcZgNzZ53
bibDzGzPLCerqz6xYePrrOOTyw43kZVCz3915gzbpw45a1FtZmbOhRvPJwUhMosTsbpeAbFqf3hq
HxpkMIcMm/LHWQ1lfwccftinBvmh/YkBY9ZSfwBCJJIEr31Y3k4aUoxAx+IyYuZo67HUb5cPSFYa
6SvdszETcpX/i5vY7dtXIAHmVtvK9QrPyNkxvqQxZg5080PLsyyY6evdHIleyDsGQ3jgG2TW/Lt0
3sKC03lxac2PQK3T7KAAOmYUUEZuEJnusLZJevwjauiKWWN5bpDlhknBA79FdQ3aP1UfT0wy/2V7
vusX/EKFTO4pVfCDWQ/57xEoxhndgvN/gHVH7j1z5Q1HEs9nL6Ok62A4p3P2KDpl9GDlC+LrlqKi
ejIuSde106f9AsEfGhOA97ZUhOyuSrnTAfDqHCamQS9CS5GcTBSyY3u/yBzRnS7j4s6aFX+7s0+z
nLPwyoVG+idvXu35WZhQVQYt+ZHL6DQF9ZiewRr9guawnWX7zdG6WRdigSvtLotje58ZoZAcslOx
TDS3oc+5NX6Jcc2ekShYVu0n0VFeAWTMft8Dbz/sLLLEnMZa302vJB6iZEKRSV4Q/mJo/xf4ykM/
QrHYywIVutoCy+us+5aaaB0pSyk4Adbisv9qMs483VSKECotXru5Hz7Kh8YaLv0RZb3yUiHuYpi/
LTXLnC0bXz0JoXerJm1CErJlL7gws36l7ROVRAPSHAOvf/Mp/W0dl61Llz+AuzkGXvKKn9zdzedy
m0vF+97EvsGRn60Zz/RuB5TDVZox7fjLJngd2Hyhrek2QFtBOJ8pAiPuwOX7LDsaPa/CszFSjozt
s+Wr34mwg7ojwsCVc7x4KDC2+TgjdUdITpU3MBPgkx2Oj7eKKGyO9DGLYTZrEq+i/aU+E0B1Q1xG
KMrX25ZTNO3d6yh0vtlDmy65wdivqwm8RuveY5wk5DJKe5cLqT1wo2lcXx96WooIcBvd7FEWzfd3
6MBkSYJqehWTKqbMqSRf69y9zFLOZJK7i4AqimP4bHFRW6+yxVl36hLDED3HVAs15cicw77kqnw/
2o0nGN5f188mz0FlbALZtipwD7KQkArdVzCRKj/P7dSArZv38vpdPB+6GGsy4Cmb+90tE3qfhFvD
30uIfDoN58OI1T1/2bo/HALjr9e/t11bKLFKH4gcovSGEnLR21SwqIl+qH5mV+D1r0BqF6aplC9A
GOP2G04oHlPznSq9t+iLCGZnhnne8THzS3e6l0CLAXmhG8DgJwWUh6+rC5D2RaeIBbuyAncdTMLL
sO3iA74wRJFEXNu1/v2kepY1VcRSzh0obrHiu3+aTRXDcgUEn6TFnaa9DZHnY1xC8R8q9lCaw27s
pk874O3YjJjv3vnSLu/oy/fbdE25j4oNGJBQRq07H/RHipNL8zAyhd8nsbAFB3T6Vm56fWbZqTpJ
Lc5OpDrBhEkiuQVS3zZhxmGpB3N6FxUM3fviYsq/8nVXDSnGmnajqP2uzaXxkbbBIE9OnTkcKYk/
X+q0KWYe1YAg4fYM1DiJsZCiN8mrcewjEnW5Qnz+VXq5/Ys4ua42U1lhoePyky1Mey9Scc4YvVcP
rsOvf7yT7OQ0IGKwMIHO5hAny6/4CZt09TZJZKbxthm+EDwRbRLJSE5YZC0fwFrCdYEKASQ0RSOL
F3I4sxv2XRpoHq+OfOAQ7MnOqulo61NOIb/M3Bl1g0JVliq+a3WpILFbkr58xykr4smouy4xQau3
0A3aMWP4g69wPpES4IH+QQtDpi6yyprKAfdgRbWIXqa+IhmLzUvYXpJpdpsOS9SH7nz3DZbZIMGS
As51CkSA5fhFVyj03lNtD6+CY/irdq5ORbZsqU9OTbO5eNP/VoZA0WbroL6eLLdbUgwKg0GP8dDR
QiUIwyFEBTq53j1afh/48z4Z2X1lp/0WtppMqvsD2ZqNrYPJeCpdGOrJlEL5GIhirWZoRu6zZArZ
oWob8jVCb2eDSoy8OyhfwoTi95EgUoareRXjxVPm7473B8CRX5iavLf08z6iB+6YbcbKXNHmcXGU
PiGvwO5lidyVjKA12QBSO+EruvpwQaP9j9CfxtWkSkXVQpNX7dcS/gULijRoGUY4C9VPfGReviTX
tX7PSI7goBHmqy5kl53Cyqcv7vUn3bKjokRne0H5nB1fGYUDP2EDyl42G7XpB2itA1vOGSzyoOpv
YGV++s6W1Wc21swJm+QRfkJHj5gaG/VZft69cFM11JjfpK/GzhaK1JDSe5YvRHJQcZAiEiIrWJha
eOX/zHBAzUJ7WMZ5NE8OT+EpehIqt7EJrqS0GbT3TjP5vQrVd1GiEriYQKqO7x6X3yzBP1iZA6l8
jLJbC2p2Iqn73kPvRiEuCWUmfh7eBgpxVvH2n7dfLosBPk1V8d7CJ+i6jywz8C0jR0NiZ5z9deVf
ZTQW15admhlqD4kciop2O9d90fWNK+60pucd38Tqsy9FI2VbJi9C0wIOKGo65503pWJ4w28MQ/70
iXaxqzzdfHIRMOxArHENtr8kEevgjvhzmY5cw+YYP+Gnt0FdeclHtbTkV48BcNkt8odANy7TjTN6
JHAg0nhsED4kMHJCWKE49xwQZCv+hE88HatFMsh8dEaGughwx6dGxZ9yMpA7bjgIIfsngcEaF98i
Q+fuqA0/3esvMLjOx4iuwfly0fnvcw4z4NxbE2CUlhixiFyj+l+6AO6TC1Mr1oATzWsKazdZwBTz
F6I93lwzfGdd1sKC5fZUv5/GurM1RyVfSY6cLUCJaQ1DDqI36A24oylu6DIiiB9JsGt3rN4YFnd7
ZfjB9TNy1g3/C6Z7IT6uOYjoCa5b/elfnrRMKqIEym/cosVeWc32RYUm5/NDL9J2WLa9Vjfz7YVM
kxguHvJvPLjeNpcAi+lOap7q+L4GlPqabi0q3Ly1yBEAhsVIYXapfy2k1dFgvT9MyHfayCecx8WV
hKFUjHdvYXUeDGffWJs0IlityMwzMX/timZ87rdOTut3N4uSpOmsfQTA4TjYySSuyOGlGLfYpcb8
hxS06KUMlTfde+tS/TzYnPI31aDzaD1tpmORTdhCOxPz+tFCXTWOjfxL78y1ORZ6xn3Q9qVzYJmc
q9syms7SsSGne9D9mFHhZGkc0JK2dVoQXd73HcrcYe4+a45kilv50xEsYR7KGWjUAaiCvKmVFffH
SHJ7tcwaHfxd+YXIkfDPHdwUgUHz7VVWkbCUGAW1ON7ho0q/9eSc64XjOda3skrCKLCVnpKGHfU9
Fc43CwefLiJdMibgWcBVCqEMqZ/59N/Y7Uyew3jxzWruf3IxlD5SLUuaJ6sUctPHdQ5bbu0U34HS
7czJ5U7LcqO87L5pWSXXNrGybnaDGFb9gInppvfyRmfuB1gvAGg+QUFU81VVwgMwb9jI+LLnpjq2
d025fuqcc2bhtUldTEk9T7Zj+qlc7eXVXUGjBplOIIfyDhX2BtMKXdQp+VxADlPeos64mN2JFz6F
ALBp+0QlIYwCLpJBM2d/sJbD23/PjjIdYjRKOtByykK71hFgr2CeRrmdSEP+wvQ3kkZwLJ5TUJa8
jg0fY0NbOTlhMOuhvDLbnuhyTgqRkLdwN8VDnoZBDUYwCIkZVk2351Z8b/F9oe8PlLsOKXB8IMOB
NLAdY3b35YriYavrihFqFdIX1d2rqRzZHLewEHbsjQ8zdiA0fMTBkFw6Q7IXQ+ycqnD3uQPjW26b
ypSeIRMxO+WQx0kKbX4F5UuIcimkoifDzohALuL6YbL7DvOEHmfqmnlatQpNKU6J4CLhG5412PnF
x7iLeMvmek04HWzDPRLdYqbz1g3VCQkv73NGZsKC3T+qMidPrXanr63xicYBwol8vOc9tyND7KUy
DmWKmaRQ1PcYopyQgA5lLo8UuzywhfO/9EeVX+wHM/ahbLvpEnQ0i9pZzELDgLvudbVxgwOREjqB
Zu3+6vsfvIRbOPs3UEwKTE6dN0NX05r9ETufYZl6A6VjHzpM8711lobM1X3GsFhbIsvSYdjs2CXc
+khxc8FnQaZIfQIg9dJRnnd5GoTnXwJ/IzVVJkfyiEUT3zOM0jI0jY7Ah1V3UXS/DBZlhsR3oUAa
+vCtEw3FScE54wUxpJ+ZJdyysE9VeHAO9VPYGhJNx0tiI0XpzSEmGfrRRIQuArt9Fn5ydG46IOJM
axtPNen2JL98Zn+KAHiMHyCWWKjS3YeQY0/F7mE3svo6nFKJjjWi8GT5F+YVoymbrI5s9QPcPhxF
8Vv/gSGI/kwzne2xz9q67TZUdt1GQvOP3AyCdcpkJjKN4ZEL5e4KaODMSP0wU8HGXe6Gpob5tq+N
WJspG5X1dByRtYPaGi7UY7AjAEyfaAWHe0qzUfTQjicaCdAm7QbThHObJpuZJM+qrDHGCnQgGJZK
yfklJ81x3WagDRRZk83KEm1q3Jg/IcUcX5znM8hmvN7iLQVD+r9KBgfcVO8dW2HJD331Y5xV0uPP
5sIWaYYynafBuFg+Qirw0qzeQc6P2SbzU1fGL2Ej5Jfj3u0wel6IV1GGWuoKcXatka5beDJ/6zw/
o3t+fplzVBlCezrWlASEN0tJFT3xohXOY0P0YJFPfcI2rhHXvZEyhwPR2czCcVlc5Bo6+9Xx4oXR
Q8XUN/Q1Bcv89aA0nbCMYcxX3+kPKYs7V+HUCNOzUpsQ7uu4d2I4uijXrozD+G49CDjIJp5H5mz9
DvFzhyphdef8CCG29CBO1YNwpE5p05B+0dSeOA9iNDOyjhLTnbrPw7R7NCGNvaiAEgiNhpaNgHVK
IabrayQkyn1LgPLN7G5DiwacAZj9uV2yQyOvz7byN7l86VZlOJSbsJk0g851UO+2Oi3hJ3qtLMs+
W32pNTJnwhasAX6GiH4orBnosrviYVBXpweWb9psi73kHjzDV/IMJuvF2ZlSHFEfWAD2fcfHM8xB
/JzJUXhKsFonZl7HVxpRAx3Xri2WZNS94v7wTzg3xkVRvVNDPn5f9hMwNIlgKsZ1CvNC3ka3N1tu
y/mYZRPBxkqgocllSzh9I/9wiAw9L7BUmlPgFUCUfAbiNrxEwyies+NBo5Ypsxrvl6Ww026HnaHY
G9fjPIT/NZlWRbOL3gBW7eQ9O4n07unfnp3u7ZQSUvTyb5igaPDn57LJ0IFDOnPNaclvKl/xeg0c
r2FggJ6kC4bJQ5n2TrgEb8376ssd+uTAj1kCdyBZ/jcP+8zX9AcZFctXInpr/IsSC1lAoHXe5U6E
sHKKsW7YOyj8UgspuUMLnOEcHO1Irx845/a5OUvyyQNQ+A1RjsRK1zbMzn0A4AGf+sbFr77Oc4/i
qNIiOMtglTAv3eEv+E8W2t1kdWVwxSZxZXqUsyVFfxC87RCYb44Htx6NBMxKB7Y8+wq+GlihzaZO
iDBnoOf747HH0KL8+hf/yqgysgP/5QuO+MWvBMoKTMoRCDkgPnnY6iJQpD7NytU7EqD+tV9zvqbF
Wo62fkUrgY+Ns7ak0S45T9vKvtcCWig4tmE4UC/mcpQzBgQ4qz60p6RgW5N/WqOBp7oxy/Ka9Izh
umWqsfmaFv7nfV+/UyPRRYPB5DjJmeRXi2tnHhaP2hYh7Ptw2a0vgCsQXfEzxj+4g+lTHTBzJNKc
+C4AEh/6FVnulVDvmd3NLB/EHqHtfZLJigwNZjEWVeeQlSshyfWe6qN04fKx/X4KD7hJH7QIFzEA
EwD7IGA7jZBPhpv/gblQTP9gtpxiz379LI6PuZidx/5Qw7sT9Lb/cfGApp491xB39cO5CGZcjLLT
kw3psthtLx07JQsSXiFCSHn2JybqqFVx2LItP+gOczZ1bnL02Gz1MkCraac1ILovqDbylADa/a5n
F8OOD74lRz5LL887gLEtXLt1sxRJZKgvKhY9PMCMSFDRyWm6WHdypADLMguQLR+bbG4liAYf9Ed3
drDVwzdG2ef20oWEqvRsXdTKN1CaR6S/b+/uUYix+Wc0Ba73KldKxDwELOZ8YHhqMXGpu6bfSOeJ
m3pJtMcI4NHILbqRvKowMZNJQAJSKwq3cy3Fd5FEBj4fr9p9FJ3dNsWZZzNptNlYsejHIM326tho
tS5vetsNKZO3gi3DROmidjJuEAVhXwp9d2dWOD2TkAek71g7/6fSMTO8moYb1Rxl9G1IeTWsjpbX
8w1UvNAAVUsoz5ri3J6NXEU5VKy1T+3uxTAPxYa1UhTcg4KYd0lOBRYFwJBBRGXTqLpR0ej7o8ER
gz+CSRh0tpO11LC8z+5gBizKzP93wbKB6n04nxSBp562AHxSPhlpJPV+kObVNLZKYCm33dMjXo8G
QrhEk9187QoRQAonijwdS5BNrrVtGKzLW+hZDD3FWkKcuMat0Xf2q9IwewRfGj+oIAbBe8OaeXQi
dHh/MX2hgDKRRTOfVkml3MezoB85MyKseN03RyqVLsdLUMHbQppSLE497y/y0XOT8xzNexkIsngJ
UcD7bYwJDDFOpzELcZT4VXNW3eWamPOduLCgQW6GG+WDg4OXg/OimzEf8kqhgvoy8ACNwV64l/EB
KVDWQiIDNivxJ/HD6tiq8KLBMQuaQrdiiWaXvY5rNJOPPKOObswfzq5dZANv3QaIgK8fgwkPYer9
5emcf4yz8dB0iBzKKDfL5wWsLmJbcFD86L5MwRcsjfU4uq+DwTYf0vWQ6QAiotrKws5AtD5j8xPX
Z3LLHOj4oMnMgqk74fdBiCgImwNpjHeqojZkcsNWEmWsFr2uuDmh7o6aGnDWrrYqfZBTWkgjU0YR
vi67ZT/1tCb9gO6IJgHkzsE2xD95FxFNI4+VWTfFg7BwTM3sxE7ELTk1K9ra7D9gvJ2jG+bhJAc4
T6slH6iI8/p/Yyymt2Oke8hEDMACp+yk18rRaXAWzgSjnPQsQTW6d4pE7CtYZjjih39NYav+S9qj
VpNMsdSQH9P2s5wathDmwy9y+kwhc7Io8DrTR0jFInumnK15/BW5dCMQKBPo9zaKYZeU9hgX5Zeo
8Bi2mn7afLp6tvLmI3POlDvHEkEReHnJAk0gzVMaSfXaUgU5Hevs2nFprvdNrs2hvqRoCArrH64V
dbdbM5Gi96zl+YqzrPPwNndPISI4iEIHS8GcbtW4pmcgMEdtY99HtDgBAz4OZwR/qzMa2XNdJdMh
BJGjeLZOg6NmbJ2gi6b7kHK7P8bJVqGViQdQAzCnsc0AETskxSZRQhuhwpxGgndLLW5d5vrDoiC2
mPjnD8u+GTQoJK83ZiuAjANzBVdhOVC5fzR1CWiKouzrBpwmLCIoWqwnwNZB/l0TY2N0okcydGNT
zwNEwNXr+THMNlWeKaN4AjckNJRJVdLaeLrea3jx1/zpdAZ8T1uZmcj8nkribyk95O3sa1jzmmvt
CMD68dP+1XatgtVoI9CnNbYQLcroRohLZmJK7DSkuEliyksi598CYU/3g5GJqAVsGTimGMciJU1T
Xuqehxn2zLn6sttXuV6oZG+XRoYReJ6mtX+yITAkHmGiWkU+np52ZLQG2vW7Vcn3w0msw8h+AKaB
KXzSHPHYuJ2yBPaZ4o0TWvDazcQUYdbmAqHcwLxGkIERWhcrGF8CbvXy3pJQCo3VTavywS8gY7zL
g8+BWvlU6+c1xcGlKP9eZQVznzscH2bYZd+Mqe/JlrT4MyGwNmZ2UUVFdY789Yqva7j8yYmr5VJ7
TeezOLXH8ZbCiloGhdmEqYjnMBLjJS9BjYGcAkTZGBZV5bPmEYBs5UHn/HkEL7qbGDgvah3XikCu
c+j/ocdP4Lx0vC6kKxDk2EEEhK8pEXdDeRnC177HZbNMvHfoFoqDcsSfw5zT7tphwubrdgeihBnX
NqZFZ1JXejJMmF2w41+EISPrWg9G53/jYvy0ewi5LsTp8PsRWaEXr2U7A/fCs/DK48qM1/p9piPQ
68KtoTZFBh0Wh1CxoJ5KxucejNJp+K6l0ZxCLT3gqFFnRwQ7Q77p/EZh3vzMZtU2UuViCTUEYSTt
O5w0Ksmjcm+eufucfJd32jNb3i3bI1zwuuprVRuf9/MLfmbYfWM4HoaYEIVfFgiA8QqSXIeSRQyw
iKz1/fRctPhsITmKGKRZWFqu0Dzs/9u3Gy0adxGv2OQXMm+CY56KO+gV43lBWYvmH3EiUiKaXVjm
vonmB5p4tITz9jFoDOvSxjCT42+Zsj2G7M/+eW7i7sXHwpsRAmZ8Xgy/ch7skYsxTt7y+7WgqONU
9knwqcgWVa+sGTuFBWmB4LMx7Qs2h9IGrSsNpIAwWDOCqqE5B4mL2UAQ/6HpDzvVwovaqtITMgN0
Gx6somI6ix/4zsSpD4R7PS1g8F218/IttddCWL5pIp+HPLRSU3gKuWLmyRWEuYg7PtGIntmujwqw
l/3K7iBX1qK3/epld1No4Gf6Wl5YiXU2mXOPLJfLEt8kCSXvc4gSp86hy6CnMWnZWsWSo0epYc4s
6EeA5qQDPXpe2gHjZ0GWAHpyFGJ8efypVOCJLp0Mv/SErLNebyPV56uWbSwAi1zkQp8DZ2MshdJs
+pldVQGFt/ZalUPW1l3+pFrBBxEcxNxvmZTw2ebeW1Pl2JWq0zoPmm/0HVCMw5bLodnTvU4thufh
SIZ6TVCJDTzaEEZGRdC5AODjetpg19DhyqTMfqIm5IJGg9KleLS6rpuOPzbl+WPESSy5p6gIKj7E
/izsvQfasrGVTfaagKYve+9ROnekpstBoHNDcVh7P6FknjoNWLuw+Bo/o4ty5JjxWiBG+DHWPdXm
QFDlGDVtgIHoCPsA0i+j/XZI0GQjnjWfvxCVJOJ8B8SY+5pyh8ImvEKDUHYJVfQ3PA4E+YQRfSxA
v4Ix14kk6BwvCmyqGr7kfdWnQli6EKuS07vqPSN8biqEduvV4pra4BI2PYOD+wWWGPxO5nndyzRs
1UVomWYdz9FSKGQOH8krEPNa0ZlFJcWQir1QWX1fxoNKzGjrpC6OHaBqIaATk3zYh5630lyvdGf/
xvQvmNYHFbLqEAZvDHI3MTDgdgVfMRK7oqvV6RhB63aAR20g4KfoKpKNeHS0dy+3xw/QpprS+NYb
lDhsjNMAXPYgjv5y0iu85QhYBy/kESJzRxdUUJvmGKJV+GJItXVeELkiKb9RpwIEjtb5Ua/7gqqF
14lwt06Gd4l1a01IkR1bACy16B3UVYXIfRfGTzcgbh21OBGhdiuld2E3/hkz6SbZlV2josRH0UU1
MI8XiC+QY9qxKWAWCGBM8TReIca3g9ZiZZFRq0BQuYabAyC1HJgg8qmh2E7KOESSoLWswAPp49bt
owlWkIuXKSxm7N+QZNxUGtUZkznoU+9fovKD6+Se6IpuKUYBbydiZO28Qo0VLgbw9CeYxl2Cw+wA
0JYGmTrFp2yJ3RFlcOqWY0eMUBfUEGVTgbjVeZrbV6pTf9sgA3oik5Mt97W6Kt/yOU9swbWFS1kh
MUPhLg7RobNYHCp+cJTM583aqZRBjRF88RUpNnUJkckkmBfU54f7h6HxAPefS0HHHagFu/2X9SDs
ozv/6fB35eFOUw6yxulMlUukggYZlU5eJpJBq/RzCkXwhoUgpByge1TaYY3gUmbPczYlMqFrdYy/
rTOLgmzvCvjMKwvKKQddplSqPaI5AY0FvWES0jfSdIcU7lVi9szcWMS4YU4isR68uvy/S9pCI1Pq
oidjcLM6e8DXnzSGO2XjScJY2URUSgOi3ndnTFnzy87W5904xlQxR8YdCuqz+nzO7mqSTmOifjhJ
I1KWP3xKgb1pAuohb7NkDH9T4ST+lNeF8k4M+nowmKzPIc8sOnp10cbo1kkVI7OwtMfnG/uQE21w
szK7R1Ux3670N6SlvqaHRmWGYgJpCwfjhR4Y7fCZkBUWfPcHT2B45jbYvNVYeD0BVG0Gl+/bp9fA
8CZuZaukX9Vz78+a5mG8akLHvlQ/dBO86Yt1xjUUhpr4ffvQj17wfWr8Cw6NnWN7nSyUcICx2UJn
6aA+safegGkeFKkBwlWE+cTTV04ZirMnbGuJZECG5youfRXG8477Z46U/jr40LVtRMHAm6heBF9e
eiWx1okU4ANuH02TNjo2SqS1qFC5XhEHGTiKwhsL+Z1zltkhxYgABHPGbQfsBYF2RraC4xUeS1Zs
alR+eSbzIYc3vjy/lCb/FCH0fiNRS9wcOgZnU//3QIn9D3/WfyyP3190FVmHs5cUAw5IgfAkFZvC
bX5Go1VmGvKPvB7/zaa8zk67b/vl3EzD8HWZvTGu/pbTQQkDI9yUAK3pKf2a+zqrgy2It0dDbSM+
ibGm+pYQRq9PnOD1LJS3xFyGcPS4jkB7fJiQNGb6XMBarXQkaQDaou8VqDREgjrt67S8MpCFo6As
h9QPWmC1tUpdPSzRYf5Sof1w7rGG6/qPOC7OZhhLXCjr2tgo46ujBAnJekRGkpdooZ2GvvPfRS8+
uCwAvSupKsWKoiGGV2jMu2FWQzuMUxJLyO5GQJSCs9LBL31PFOCkS0f3nbdX7Ap0fQ9yjYvUsoMw
jbdhy0xC4WhAEaNjOrYIGrVzyvOyky1qnj/0e/9Jl3+Lxn+lUNCFP4SMF7p0TkMqZ64/EPZB1nNQ
GkpLY41Lmoje5G1iqk/QJ+a0MYAC5mNXtdJUpWKxECiR9ssh42dQoFgqSwHR3N30gxjGs6ZwjrTI
y7LEq8q/B7TRQkI7Pw+VC/3nM4mq8LwF724b/p3Y/Rt3ADOHBK6/tbWjbr5mN6iDfaBqPOHonIw1
JvMgDnFunquRuQziMxeob6ItyJ+QtQNXafQiP335+qFyFHDtrTDMU81ryxSmZJaWsbgZlktc2ciC
+qbvUsUXSDTuuIVdN4i5jKLz8RyMp6PTOfbNsV6T9nmE6BuM6NrEdpLZ09ry62LXJiAIgPSvkga5
NDXFifZeMTFtdYbXupze5r/DxC/NcemDWfoEpXmC3wiTHrTfQbNlqJ1p7nTJqx5gcALVdf1IVlIT
ppvx/CNLNUEc2QdXDDPHQtoQ1FJALGxvSt2wHOn6vwRWemBlHVdKo2qc7NjFLsR4Lhm3mzIL+Etx
0xusMSWweN2AE3VeZCPak4bD5zjJ7RCYkUUXCfCR33AixHq7Pm14QhRSc/jyY7HodlsEWOJAbdLT
Z75INYyoIVpkrxcx0toa6tiOGsxzRImuvPRC43E+wRpHB5XuP0pXeq18DkFpbyI8bjLdpLndwpw6
bLBqgDvhXCnxgM9T2ZTH65EDguSr4prVJe0kYJewPchLxZkkLWI6lILW1jHwobUb2NQoOIoNNZdB
2lvr1msnd0tC0ajj0QZHM7bZrWSIrFqFTP1Sg3FW/O1upJ8Eclf2buEQ1kqSOgrcxNrnyp5PX2P4
yyLryj/YHxHgF6BmCCsuJbO6Sk/CeNItbDhYEX9Z6fSU8NlAV+lngxy1yo25zLG2fPeYPKIbIQTt
LTT/stkoz/5nJgSTRm5nl6AlRlL1GLD27fjJmZHUxwuih2Qs/Sr2ahaOckg38O+wO5cYDlb888kV
JG6acJUX3sfvr2sF1PMj5zfSgxvnYjomhkLCq2fZ5TeZwkZz6h/3tP6JgPWkXxHV4uNfPp0mTapP
bfAlx/6WZqckO9R1ftnFj4mrq+9NRjdhf3Y9hEehkcJAtuWHb76DO8cjp1zErLWK2ocYF5W4Pq1g
kOJOM6PADdukdtI3Jp8wUembkoSqF9PdHw67izfi2L7ohCo+3thr29QofISeMJcr6rTQOwxGM3JV
WpLbeB7xwXMaV0EU8YnUAeW7hh9T4dR+DzBhRY+8OuyyQ+2NOlBwENO9bobH38Gt6khZoRmxehBk
UuFF5uPaPoaPeQPL+UNNPnFp/Nvos3LNRiUUSVu0AIwU85KPGVNvV5BCsUcmz1l+UUgn9lKWw4rS
HAZX2cPfnLmVJ265AauKae6NsGooWXrDGWLQZBWt3Wy9QJOwv7bS7cHairPHHzMz9JDdlxt705JW
APHzCp9go8Hsx5ixvupgCfTSZ+qbPtcBRMbvXNVm6EGVDpBLmv0mGmRgbP+nU2tpCPGabZrtBZNX
44SGuvIjjMPiy27Bea9Rj2m95BLmqCjpR7kqlfEGivcJJEXf3RqcgXcndpgukTdjwOPhR3MU8b2T
qWH6BIzwrc6LQoitTlbvUuvrGtSZ5K95zLJA8d5cBICSBaSdjNWyOh7CDdOIZ204MUgihUiu6Av/
gTIeTPPxR5ZdFsYiOPxbS45hOZ+TkuruzgA8E+w/j8ZQmPCCHw2+BzfVxFk3Tvl+Bk/aCfG0PTzd
t5rMtlV8Lcksu2qlcbpn31pz9TaU3cRKRJ7p3Q64FVxh56/AibRHmG6afCoEKB/FJMTeoExkq1wH
mndJmms+CFWyM/OLbGHcQ+iqZzWPkcaukEQ2eJrsYWM0IehUGJ+3YpERoIEShtmBz7IPB+Fn2FNU
9A6CuImw1bLCWlcLN01KVPrMFSg8AIoJbgYPG8mJXM+kBM8wmkLgj7ZqW//e5VBV2RGdgTwjlUPZ
BOkPtTk5f8PNl+y+GtMe/tJmDs1M3WoaDrwOIgScdMtxzzCvWKbvJb2s2pfJqOqcDLWaqzt5qHpR
Rq1xPpgVqy5+qXrHHIGwRq3gUQ2uBYXVPzvXmWPAvq9J2jnTu7hmEUo3LYWbb5Et84jCXUUoEhjr
p1zIb+K1qfj9ffWqPX8EZ2MF+8LZl9D/kCuKSrmwE7inH/UgZBFsTCzMmlnJCDBApS6/j6DVhS6/
ACL41owHWvDwCSdrNPaWB4EtYoACBY0IBqgp3VMnsrQkPKK1FWOtuYjgKa1Eap3QGBwzNuENK0CE
kAb3Eh1L6AGUO9CrLfFTwWRhB5lv1vTfgwF1fsyeGdZKeh5EBtkC+04nBnZpHviS4kWzVq4HYDU0
O6kmpNVhVhsa1B6xVXPg7zUWw5/vBUUX4u6QaUKGeulszoj8DjfLR+2SPGhfdr1SB08ufO2kTYpp
Kgnfwmo1x8I8ew/KU6r6oPGGX1GQcCa2Vjk0bs4MyvZ/mDr5RBdtLbvabS5KKhoZ9kidI5LQDlRA
E1dZI9bVgwoVFpQP5dluevzyqox3mou4tMF48TooClyvMq9XHfrRjIuECgSbWDndHVltdjwreMNM
uFRe9Ubl6zvTNxZwE6yf8iizeZJSNGNRFMqHneKZhHKd1s74IakeEWrzGWBYmCpT5+5L6uD6H99e
38AMdHg6b5KDPsZqZmkkKm4YGS2LxRLidBBv5k1ubOOYcMfnbCPG1dolhav6MudJ5gensl8Wjkod
rBsducaEFzcsA8QMw9tmH1UhBb40izqGhI2deN6p+Cb4tS4jRSM5gFdR2PGS9xSTyqgwooXM9s4G
Fk/o+hJC19P2BCty+cTNvfu9wkKN/L5aVIYuRdKIf04s8Q/3DfpqGTZyNJ7D5nf/sEXeOOUJ9hPr
sv31RsEHKkJ/uszAwebBmt65X03G/xPz08Z19vTtPWhKqpt7GpFJQGUiJ0AfhAM58vQhM5glvnde
nx0f3wTrpuv2DnAmqsKXCfllrtC1SHZaL/xD/H6uDjAStVFH1olYdLa8kRSR3EUygujVDcyqELTh
+VamwSguGhU0AYFmEapweHnIC9krEnbG5Ut0zsVJpclYF2/x0hnWyl3RL6ZDhQR0mL/epIWwC18v
Nbrc3HFjuSdm+whl/y1kiz513ovs7lK41WYACL36ORUpy2P+6a70pWd4+ttZRlAyhDUD+6uToNe+
wRegGqdzvApyBMSJuvvfdImQW8HfmbD3+agUI4lJxj1Eja/V1wfaUt2uthxse1ufrWtvpwzBzPvK
POlcFzDuZ7IQih6+KQKgoqaotI+je/HUr4MZdujYNxC1zY1Fgr5o+XVnpSIhRBK+N3juX0AB6pR5
MtWX9T1ig3MaG9Z24MSVQDCmG0LAozuLpFKU7L9Y8JBhPeIwgzsxTJNWkLXPGMAtcXSt77vFVxFR
vknj41rTZ466mtcQaw2xD+MJhaOQLol8IYDVQCXlBWinI75SsJYJWDETVRstW2N+I0b65dUnJ/nV
EmtPCYC7WYydn4dxAlFHScRIu6pzewVmRX/XUVjebo7+aW0q4NRPdjcz3KvOXh3GSyaSaBJTGpqJ
Cw7Vy4/HznVvNiTxbT3vt/iZaAlnsV0Ny4oPBdn2uwmsmZayZmuECUf4XvOKlIadVN9BetZ9/wTS
YQf21UYoTf7sDZQ4bsFmncbwP0+WoZY/O6XNFehxDpwezpMYFoWPeFxv+1Qw7wKP+XtVYu2MeiaE
3Wtgipe5H9o/Bl0aBOEtzr9RjXIPg8451qkUzjTUeus0nTdeFu6hstTLs5S8OMwgj3IdvZTbhZ8A
+BK22F3Nv1wj5rOwHxALm5XW8biZTKl/bo1ASV6FVocuYOoRyiNSbGSGXBWPfVF5cxkLhfmX8XRO
7ujpm2Qaz0xvhgqgh7zygkU4mUr0uvKlqury7t2YOmHmj6abKJZAgT55VIDnu7fwSbg1Utja7IoA
WpUgHn5iqi0U0AIFgVhxRQI0sdd7Af9NJBaQBaMDGVXeV5DyYFTNxEQv78HJNDNp59hAqSamGkxl
nB5I996VhjBhu7AQJp3DE46gyurcoK41ePwh1PXbqVvLpQtetWw1JqcmEx5q0X+YsaYAERzeyzFr
ahbBj+t5ZVvhvuSrzm2I+4r8qr+Bs50llHJhnRMNYnkkNtMkvSZjxuIP27WpyB7yZC/oASFxuwuQ
jmCEn+g7M+y62qbqlC7iiF/7KNM4hmmH6d450SkdRehWsX+BukdPNiR/iPA5v1R6DdHM22B1GdH2
QpfAuGzZSV+EveFU7lmXwVT4Vi+r34K1W6Cc3AZTr3/8ShsClG55G37H7ZGqAfI0XM1MMZAbz8Ic
8lWuIlAlVv2vW3LczEhMjqs4QNO29kJPC5G3AtU9a1UHt437qmWvkN9BPr62QK6/FmHd5OlbO6ui
pGf4EY0kI1AQzj6rKQyi3XoueQV2fiVFNAfQKHpVOFZYGNmTsoS0c4Zz798arOpzv7TOByAoUbi3
D7FkOWalGqMefle2OE+PRjbkKj/chuLczKnTBmteq2dr8E6ogXokE+bR1knQp1jj1rquZxv28dIt
+h8G/uLFbviDligrin+4ShGYNOYNV5Cm1r+gm5YwU9MLlJUNPIQw/NjMFq1vbp84+uSCOW/kQ+zW
XA/J8o33Mm8J2QeBQ7gdAtPXSWkF0+4TtBvdyaomPqDoVoVreH1pG3tQPKgdd3633rLVH1iTKkZN
yVtQkAEBkmjUtvY60/CqlJZJOZbHhUq7A3rYOmYzPGuzlQia0gpjK2HemUemKv9xmOMYgUxQNnUt
Q6e1aYmHN3RaQ92o+cqS2/pmVA4CHCXwzUh75u7DrVf/oeMee/4jlkNInWPxI+17IzRkBsQW3j+5
zu33SMUkslYL/Ce+L8oJuN9NK0yXnlUv5LLvkzSoEv51fcjmZCqG9Y0dADKwWRcRIFZuZbCNtYXy
vCFpLxE2MUmqTPqkwGzPcINYo+RP6LUzKwZp7RQwTeh4tyykka7T8u7UssAGsG+amGXZzNsgMYq/
M6XSgmjmaGv9IC8zVftHJ0Zhp0AXcQ08pPx6HU05rtaNPRXgz1hI0JgDbcK6TlAo84SB8WJ7/Xk1
re23mo7Ocebi0TMSAqE5m8lv009ZkbKSG2V28VFKkGbPwU34T0W2XOhR35qGB8KMKnuZ3h5yGGdZ
C5Thamh32tm/pRFFsJEXkqKKLRD5Up1cPKsxTRlcTukWvz0HCMLyyHYKukKN5PGPhNcQeljJ6DTf
F0fhpM3ltry3reOs4fnRt4kgQ96vkqNojH1u5XZPanEF/N1l2EfK6hcLekX87XXbnEBBcAUbyuM9
8YKacKZ1DcglkwZddtv4GCauQmxWeAhNmnqczlh59DMpnwrZKGGDvGNrNY+C9sP2DuIy2qMm39RN
fIHucNN2dw7I/pGZWG7AXaL1aho7S7HzrKJppB74aG8ANh23KoPtWJVp0MsUuUnFx7C+38u76ejk
oEDN/6f3MnP5hvk6cXJsKDwiHzSSJe/zxF8DGXhEvssmSVtmGpGcVUb2lPTYFLYBtAY6UG/TspTt
Q/FU3AJhr4tCShh7KDJHR7EG23JTqV4ZMffLWorivhZZK+4Kg5yiZHoPGQRfm+zmEghM86MJFKQb
FixfwopbzV/DW/f8cR97sWB4NcKua6hBlaV7qhghBXs0gvl45sh0mQ39ZGFJ6I3AnKfAqKSEzvMM
gDlcfyLR+1Gcu331A4VV7Hlq4GpaSOVNsmW76PWIhypZiRbleagmStSQCQbKTy8tMZZDMlr2+FFS
H/c25z0T86CVERPZ4Z72bzjFaXjwS0doLJB6qzEH00kqBsxRzU1MfbHRcLceYquczE6V9jpLq1dz
4sqsV2nlhmIOz4g5LhDz3UCrC7pa/3DXOrWuUtRIAbNEEnu3HdDLGCmkjzN46BSigOUqHOFvHSSq
XkUH0uv6A4jqAxNovSSHZeZ+XQtWmQ+JQdjK1tTeDOdvMZcSdronXyrjF3lZ13+t6ygOqchfa+2c
nq0BJ7+hbud4f2cJAfHGWeIuU1cB3k4KOLUA55FhGgLtx2vvA1Z/Uk9hXSULISkkJtar/x6aTN6D
upWQ4xnNuO/qinZ6t7STlnp6QZrE5GbRoymXTBvSni875Jc+7OWynhlqZ5Ail3155NSxTk9TnaNo
oiyzloP9z842rMGFymPp7vNvVR5+b25UbAbqollDNMRmxwr+cg7iiNath2zyPdT9m7oyU4Dn0uSn
iFz1lSj3aFhGwYaOU+Tw28v/Jq4TLuad1QzmnpKZQyVHGQepty1xofrh4LQz2KKjT0ws0FY9Nnym
wKqLWGGa4W/eMzz/RoOLC0YP5Dr0XwjluQpQWC9JIqsweGFqOq70c+aMImDIM0cKT6hCnh6R0f3J
oYhdL/RwIBGaDhg9RKWrAextviCjTjPGfp2d/4R5b5sp1eC07Jx/NngPJkLPBgCikonQpuSXTC8+
PjTHPeXlnYuHf4Xo8PNwyeqQXtCS4GAfUNTPz+aW8HcXISQAHfNWmzwgHfXZOkctRtaBkhdTjKic
KXOxZpzZS6aph3DqBlFehw/CH8fsw3YJi3/8xzFtkxVRZNbNeISpjGFv3SG+GIKa/1ibifTL6fSG
zSqua/zXelnQTWy9XeC500RQjIhXyRg3rhzxboIgyh6FAfWQ+Rp17YN3JgTxKUX3b9Cd27+7E4wg
d7179H2DmT+761PhqtJ0of8+LvwAOqnSb+Gi0B4I4H2zZ/PsDTjLomPpPxGiyHBMo4tyCn7PDNNF
U+huZvcbfV031F+M/P5IJJThYenArzES+l5pI4Xkt2vUX76SpBMdYxmpBaN/nPX8y46AAsLUHpNt
Dgp75YWnTXUoJyNqOPLXp7M7Kd+vBcJs/R9+9w9UldUCIuoUXzxae4YIU1OuVObecRV+hvy/g60h
cOlduBZ225QvKyvUVGFGeL5WePdn7mO+xecbYRa5mqMnZdXUPku+DkAjdqdcoySF5xoJqrT5dn+R
O0Ail7w2TzoLzpXvywHJmKG7dkEGQeear6Pp938Adrbc8B0dUMus5PdJDwVqWXkNiMUgfqMDLwHz
FJ/hImsfWAFGZ44nhGv6dPfBsDzoWAUkbWwJCmesulGJVD3IHONLmJnbQvsvGGpy/bR5OoxCabjn
0PI0m5tTeYqyT/CetEj1jNKd0o591nvuxhciZ3H8CV3G869533Ir7wNUHEzwirloKOXw4DmfnlHg
QNj9m5SnwqN6A7fXVhAQwzIyotg2aECswoc648a0rylf49CQYwrnpEw+IOAZgJFbNDS6BAUmTCTW
Te0/UWEYwz3cpjvdyr5zVT5IBvJ/ZPfQ5595ti9Ax45YK5K4uenx0rrgVsn12ZfKDquR1i3oK3Lc
pKvBN5pOptCq0VvPACb/bEpAMPEXa6tbF85WZOH2dhoRCFCulqhDeDgxHgPwZWrliF1rLyDp0gz4
7TNL1Fx0zWxEBftIUXjamvlxSd+qzsU9gf+BNa2TaBFPZUMllgfnpUxU46sGAKeiF/9iRarP2PQG
Plyy2BMbshdiZDdvE701ybPBucyBl7+68nesS7KRGiCrSEi7F2W5A16oDNy+9eVnfAiSCuHt2L/5
L+gxJKvf3uW8e15pkTh4vKJb2s0XgOtTSQo1MorTb19Thq8bDqNgeFW3HwW4/FP00yu71EtxwqqC
p40eKmm4vSSA4rh5pKxk/cAgcPWd6TrcOfYVzNP0yIDmagma9h3bmf+UlYeu4Nml0asykr50IHEy
UCYj3uXm/Y2jBi9Zg/0nZ0usjADJ57jrLK7CFVuIfMuFBjm3Z7+TVdOJ2KmWuaX+pYCmDJnttjkc
HgAfKix2PU9v7XSrDwfv3ggv4TuuVGwMpj2Kcvajzaz+HaPW8PWogLZcbTg+WsexX/pAXIxjD/BJ
R4zUIc6MSTJOS5+/DpKSRJ9d8QLJ9yk3lk06JlVgqTMIXP6qGYGlouRuSv7JUYUcC1m9HcagCQBi
UYqq5js8ZNs8g3FlmPXyLwmUMSJceCgurtGv9VLf2YU1ED+uVg99dJjNTKFuhySHb3h7B3lpkhaE
nmgunUSfR3PMz1vruiN3j6b3GKkiGZbb8U/p62MG1fHzdTkyFlFqxPyVDzHWwbcDRZ83+Sz8+vyz
vAX4lzV9qAC+SCfh4UZ++L6KbEeMmNS7z1+jUN335SHBTZb9LqT9D7W2NzRZVfqcJOSA5UTVbLzB
kMpFS5LuHShsVHVFK7YebXbrx7bW19+5XKHjOTIMInRRpTfr10g6o7I7v4lprSyHt7jpm2d5rB7d
a7hYENCoV2SAD7pJmt7Dfzq6I363LaBk5J1EcVB+GFcHhfeXiBhLZqBFhrEZ6Np2M/qYKJyOQrfs
8xHTkwY3ll8TFLGt7+Q/CIcyR5/Cs7IIjvXBvtfjy3x9Tgha0a0LP2uDQ2HepLrdHroaxcdkCaT8
qknGY3WbCo83ZQ+MebVtzJe4OPYd7sKcCuBV0+s2WAZeSkUwEWJtyQoL6xrkpWeYcKDOvTymNvAD
0GFehRUW0XwLmtsp3nD5HaK1MM5jA2kFa4lnFot2WGiYWKkkwzLfSvmNrJLE0EyWM+iLD4K0FCgc
RFkdJH5m8doh85F5+iNNnYa3KkLg7GhHYtMqsCAV0a5vxeXe6aVvZqFPZulOtaWb977pdjOlZxn0
PK3fY60UfHaa6SYf/GCPdes1KXQLPZFP5g8RcsyUjBjwW1jtouzLqI/JDIJcNf4Z9IgdYqegeP0T
BEczbES1XFnciTUx3QsfoKBVA3nxWcbhcN1AjQp1dWU4MQcku3oX2AgMqtNmp06GwDMzDTEJNSWa
kXiqtJhM8M37ypkbdl+CdN3cjvLsnixn3pweV4lz5oxwUiD03A2ppS0mQvD08eB7IPVxWSIWwmUG
5MgwC6H/vlXAx9jPsnuP7s/OAQl+GOsTN4M5HKazSjNnBJ42RVSL7biu8chkJQzXubZIzWqUnpqx
4q6QmRQxW0heZZILEbCYR2UEafEflxwDJubzBFLw5k46b+1+l0TGY7hLy0ECUJ+aqIrYW9g4C9uh
+iC31/2EWxohxXKStQfeBfRQsAj702gtORXYhk0igEC3dgWwzUVa5EyUeaV5B6DzxU4h1B/qFT8P
FnMZ3LdQxvLMWd5DxF99YOFcimVDLD3EENfCOC4+I8XQgR2tazCuSVXBttW9f7qk3xafor0QDffk
ZMAgCh2C4rnL7wfQB88BTdK2l3QHMSCoW+L7GfWO2J+iNe2ERa+OYFOlYzuhNF/KYf3X1hU+jsoR
IGJa/N1jYQzaEswuAU9eEOVPphWiMOjaF3FTjeXUWc0Ki+CDDpEC6e8XzJ6gocuSFDI3pbGzNjf/
R6OR83GJbSoPSk9S6kcy4RBA/LhuPIIl1rXl5cJAiuiA8AYgvOF1PPVkBsURJ1PVgF0eINwYkkHW
AUiBU6BHduS00VuOgpBqfnAt5lEjNcUiwBS3H1Zb0O7SGUadGGC0nPN45v95/Db1k8vbJ1BYkJlo
NwswPDJwY/e+uaUifvicCHk8Xw1vn0TW6sR/kJz/wmzzAgrMsPDZsUFCGjmUW0sJe9UurlKjo+CQ
SS60Xf3O97QAg/8868ICO9ZrRSYqx79xURPZv7YQINuPhjOkQ6wNhzRNp4NfJVf7piWReG33XRwq
st0WZowp8RWbLj8PjrpiULxegpvz26it72x5TXqAVUaotb2td6ORub8mWwRVmEm6uP8ShtUdANt+
/Jx872R5H3Uuek3/Joi5xczrDV4Nt+VtVfVP+2a/8PoXUHfUhmNDP3i0qWvGFIFa7smco47fcDsN
GzUJZJzyNPpgxXsoVF2MQYru8yPGAs7GTQzG305pQOMeN/4Wxnem5TiHFdAE+zsOGUZ8HCnk+JHS
rCrPLn0o6s47Fe+luKmRoi3chJYMvU4Qgnl/MffzNmV1BUrFAtPDYVdbHU0mPb/bVi6wH97W3yw1
knEScLbCj4inYZl1wTc5BhhBatnN/SBljD3oFQLsi0a+dp3A/Ve7QSI1pgSHJEGgX7stjhnJpfDg
rD0pr/bHiDp9X+NwKbW3hptvA+CRDwNL8/KtmGpMi5u2SrWRG7nbTT3onC5L2grmBEGEfoF/Kh75
0nz9DpBBxIDLpOP9BoYvglE6GuflHOva4Say6yVZjW6hlsY14dfXfYgtr2BBtT7u2XAf7OZVa+LN
PDcW+A3wyxWVicfsGahDu5rxna1C43rK55MiiaaSD9ur2A3GEKVBYZ9GwASZ6BoywVPf2JNbWzUy
RsPN0gYdZ5zkJ9n7GrldiC+EXzYTL0kQBm89/IWai/t0knGK1is1tufRwbTcwWRsylGAF/VfxQxY
tPs4AqI8evuL7Vn1WqHsFBdCjiDRlwYd9jSzhEvfZgys/Vn/ok1VNa4KQFkrayZpJeMoMbzrwWOu
kgw5Es9HKpdCz8MIc8rlCFXY5lDdgr1S+TE4qrmHjNTi+PmP7BlmzYm3qVmBsSPNlK7ennZxvzq4
dVe0y1RKtGGT3MiSf7KoIOb217GsJz+U6ermoWCZteXcjO7tOPoCCxRwWFaPaOmE2upFchvhR7Yd
sY3ZXPW5ejxzwuormiaM7tRG2Qc7jBOJk3L1dYvHudGQbWvcR6myHV4daXTWykJPV2vv3i5FSotA
sX5WlivT/OguOm+fMMo80ce7Hpr4KloFy8FPFXvjP7msVc3UeRr3gt/d4Ijl/7mSTWCak54pRLUb
ICV3UtuzRk/xbWRz8yQXADx6EU3oOgAqQj+jskWyE+fm13q1XwNGnob/hQGEPhWQKYGkC9rI0dty
Ztr8E69RnRdfJQMWyOYiHFeCWZV6iFrqFGALMoDN6Rn3QBs7T1+13tSvNnluKFdNeY/dOUKiZ4zR
csEMJ90Sdz75W/CTWGuWVY8jLI3x03ziP/TfJLlxKFMy7l4Q2wQcko665lHBFvtODr4h36TdPNLk
kKwUFHsbIS/JHXIukm9M49gkqcsAHnIFdcNYcUsf4SaTOloBJdPDr4wPZ+u/ZIRVgjOD1XBxabZS
8IaKTKtdjBCokE21kGsKB0JraIpiQoS8olcsSnA7NsxieMY80vat0ALQEiN2Ri6lDuFjmUq1uEc8
Hv+u+G60X0YNrzMi9T7xKks0T5/z99EMGddk0eSEEt8S/C3ifRlix9QjlLhIweMzM6NHNlSWn+Xc
jYUwjqgIhGaRWTPTtwtGM4JQUt5WAhCyYe2WnvDIn529hLoTg7uEYGoUAk6By88l9V3lEDtGelA1
6OlRf9cj3rEl1JzuhXp7l8brKAf6AqYMEhO3rgRz2gZODbY3NsBijnOsuIL5TeJwIL0Nv9lYCqkN
6yoiTybGs7Q8j4jTN5Lq40fO5Mu7pDpoxscXN0puSMUtccWzqBKMYwdi4O/hQER0parFdI2vMiFN
73xbKUnbbNpL52S0+ahbGhZG36dWKxNGlfC4jRqX1alBHgEzkbmWueKXPjG7y8NvEM5WnRvEAfD1
MlHqZKpvtNBfle2ZERBYDy5mQQ45RDeTSpDUXlTVhlBDZenHBO24xOkE/r2iRpbZy+FOEjiVH4yV
xI7M8wGg/53IJgjNVGFhTiryd2zqZcRUBhmS3tr+QCOPknuW/XLl5JUT+QDRdG1Y1PtOHETkZgIC
SVUuSEtkas3f75R8AKzD1S40HbOJYMVgMPT94BakTGdAjO5UTPsii76NkrOcNy4+oDLcUmPI539p
ScJkKFzJM+q/v+tf2GuSXgJ03MO6sDdEbRVOn+hO7sRJb/Qj/Lbd775fSn+yVoIqXCEhI8K5ysgM
zzptYQdUqC6pio1+M/BtOqomkLP1sdy7KAp6qgIpkDaag3/wEZlVorg+cjh9IbG/GaYbCjAu81+g
952f+Z26Ao1R6XjCcLvjUw4NnuQry1la4p+FBeil9dEmwSpHol114YQpMzu9JaZyNwIl/8MHEzZ3
x4wMM5NRwYKOviQ5uXDyLjbQRmaH9vrNmFaYwVZ7ej2QBNHenB7amQxBIKXXNNqUQMDVnqo/NO1E
r6F6keH0eHqGB40fxZIJDuzsc/80g4Sp0QVeao+hDhFd3/COUJK8OmWJ9bCl77mDAVkWnMEWa509
sv8ALMk2mzSueqir4Ha4qdLSZgyPsTHM2cclmI7PQwEeUwxkW6kz9EZZBZ7z/Txg50z9K7p7P23o
3m6FOtB0XwlRNpI+d9oBxR7VYI3DiwyhHKYr1sOd2FN5G0zlIVUYSJMExyIB15IurL9kBFIeIrB6
Isn8BN6oy9YsS1DTgtzSlnKvZvLFhuaAfHUITpv6FPS/TcXy5PwVSMoBm9NtDzqlzO9T0qwxM3FL
9Bf+j1HJrLGTWtTCJEPv2TtBi9bFdu+ILrjB6Wr0yD0ReycAiJllIhQeXOnp3ex7DBv2rqYpa9fk
eSJIgL+AMPGGhaHjh5/I8goYU7lkKfybUJa0aYYxsDk/4D2EzP5Pxjb0HuJJrdbhz2rM/vLdRv/7
M8jVLyyZY49PSoRTKYdN/Kfe+OhL+9VpSFuSeuwxKNHKjvACXWyARYyZz8uLXq7r5rPZhhX9T/oQ
hU8BQ7XNas7wzqsQa2fzj6gJRs2MiFL8nYtSS0zqYrv9bqTnCAJJ61VCLHPMT6lQhjNzvKiVrriH
2tMeMdb8I9OD6xBcxFrrKQ0dFdIgZY+wVRjoLxOQ+VJXENLfZG9/BM1JeMEcZ5WA1cb++wcxs7Mr
8YJpFvkQ+qMGtQkRXejNiJXsFxJ6oyLOsI28Qdh9u2zxUmwNcdoMIoMazeyhpXrz9MOpN2FA8k4N
omu7ORE1cTZ3gnPebw5p+Mem+z7H/CYe8nJnhyYaus0NDXTt62GdzOGCWR57431lBAYf/+Y7bYQt
+NUWBhcJc/0ui/q2QEc4UoyPpY2o2NZ57jeCmkU0ycaWXzT6RL1bcpqY3+FCkWtEX3XdIEw/9LN2
9GCSAmBrMI+sqP/K1c18zhfhXGwdfXN03Bd4nUVJ+wX6QmyucVTslKmJ3VKrAyaEXq4HDIA1Nzje
JykYQnCdu/IAte3elE+FZp3/VMqvYu9YPFOik6XSKXLhxU1kFlGnixF1eApEA1lpQXqeGAtCqQSR
f6THjxMg/fNP9zanzrHKs52FyewZ1ba1EgJKVEevZD3KtjQBUPvbVelMBKuHfH7MFdggXH5k0TVa
znyUJIQnMyMD887KiDvo6zcStTEHmOicd4Gko3AJ5dooERx6CA+rnzrlr3ILMYQkCPA6NRuqHwW7
ZsNcRp65c5XDTdRdyfwHn3EIbKya+sNUFE0VF3z2Q6ZWiPcsnx4QJS+BVnNeDgKNeobrFxY1qlBI
qhBBQcbN0bJBWTh5uJEj+qD+dNoQFlmlnHiVosDeP2UON6wkuqWvfE0mLZUFjh+jlCK61KD53nK8
CwjdrhDHj8NYhrjl20w7fAE0F7jJQhLTPNyiQw/k/OgTrgMabT7SbF4HLtZxQ1K/srdTrW31rq1D
0ua4U0W2nG87erGS4RDwYyRtPEwOKZRR859Mv9ezaxcgAl3kagC4/DmrjsBPpfByhZRpS/V95vfR
E/LVfkps0+YQviPR2DweHFwloVEGrAeK9TrKw2NMbnLm7MfDnctTbY6ORM6Fz/vr/aIZ3cFRXzTm
DfvJzXb3FLvKZmBofgmSdywZOa2k/CixnGMVFj05IFsOhPnrWVNpNwwNE+NGhHCUvdveQLAa1bGW
Kae9ZG3wpEIsdLIMqPAHVcyAz7b3cTsZfDddtKRXFiLlF0jImIgsK9vT4IOC14lP6Yz7KSbGXOqb
QO8o7M9aYAQxgZ9TlejrNah8lBfSWL+6u2+RLLUJAXR4TipzIBUBiW6pDfGNUvrFTu/vSetQ6rf5
0aJooHsvOzFEdQ4UicNKI8pXKzo4gx7SP2P/9RrQkDl673g0hV1fpr1QAo9egSJV0XGS2lDzKbf8
C/Eb4Qecvd2+XTIZFdn1GQnwIxovoMkhUuKulzg27B8SdgmqJrQ0tUXFakY6XnQzdvR1t54yR1Qi
k9vJ9vAmQiSlmhO3b/wMaipwoaFzUsJJWu9MMXJoStptu6oSwa8U4UIVJpYlKUHQjhUwOgvidEsf
QcH0W4YMEOCW9jytCnvimNn5yNf7zoFDZUVfdTOwjR5A+oF3coIKkSOdUZofiIhj+jL4MJlajO7O
UfYBbte9on4RZYn7ZLCZIExrBGqHpoT2peOBgLBAE3/UTKmc2MZpoPoXhOnBjEJxLrorJRicxgNC
oNDQo6pXEQwma5ePlgSJNd+M0RkMsO617dXe4RF5tgx3I7JpzJi5+YwwtwIZb8dEtXpc6nH0jWwA
1XOrqBMdfPiIKpRGZ1rHSJ+IFM+hX4y4+94pmCAWEIoOoH6yudfOHUULmYfyz5H7fJC4j/LlWDKd
YETu1OR5eeEa1R7sSbhMu7UiH815l0alRWZCas1XH38b40Uh3wvfP5fFJ4yHpXF5XcJ0KWeUw9kL
ZFPAyehSBADmebANfXZsJa7ooXwJvDGNZllKpNrCMhH4BllXIEpMB3gzy+uJiUXPbigoLgcevwF+
mwG5gJW4ViLB+xONzU0ldDsk93EoUdnNOH2DizJp+xwU5jTiWhGQfKR+6r1BSU6jNBKAIA9lJ5IC
aQqQQd+jai9T9WLuPWpBJVAyni4eL6P2Afv+ZD4Tnyfc5M6KJqAQbYYh48CIRJGE771e7+iAhLtE
/mCC9KWEeCOfJDCoshpI4BGitYp0hKYLv4pHmIu4Dz84w94mv+qk9e+tpv1t/lqllyiTMwxAjv2i
qXOn2kUKh3Lyznt7RzixRVPA7Kz3CI0+1fmWafStGtEmVorcUdCTS77f1A5l+8Ia65e4AtB5fsJP
dFUtvjdf8PfMhPK9CKadOWTqASkOHZfMpPc9yaIAbIVwXJ6RvCi0RnWOoRQJWGCid6UaQK0K0Zi9
W8KbyF0ccFunVDXIAy9Y/OsoTrVDNnGljyhjMzwvQ+gj0E3BRY3QpG1hz4WyznlWhfrc367kftxk
eWy8KiC1APXd0b9Rf6xGlndPAe/TZQ4SOlsOhq5j3r7ba/y6WC3pvTk1Owa94Li4PYauOxKb60yU
fm1+FfesG8q5g9yE/Zu2/n6sEO8/TYxiOF9OhAEdX5E6kJiYiX1TNoN1bD2WkNamS155E6hQvzko
ygdgZBvNjx0kzhIBom0ZyGDgKPzUCSW68V9FCxHwNB7kRYaQClgHFjhV5DgncA2OqvZfbFzImslX
gdUEN1LW/OPSj8dqnh95/WaJk21lo6klmtBKfAIzqzhFhq8nLAvac0hQHUWIvsjr8RuVaQR+vzp8
I6cxzJjtmcYYQFHvdddg29bGQ9T6reX+MjzQbJtKXlTiYfYphOtDpQheHVvnL9AmBMXAwzaMhnz+
2oRMBmE2S8nvBOkJ1PBfpyfcddJX70ZaKXPclva2llT8tvHohLxzyWOBB2l5ZxM+LDnY1kpii8/Y
5vG0N18p9pK2NHSx9IUgo1EC772sZPzRFql6IV4i6r2D2HaWHqa2SKibs6Tzfc6KO7lNbLDsuRX/
VbtVKBnlwcStHhxV/ooY/dvkB5W0ZCwBJIc8X0bLDzkZYIDUDcMEHQ3LuIvRq2PnkjdWh2o486fl
etcY3Yba/YwBc91Feyu0/uKHeID/uY8qVUCGl9zkE5wRuR8lr6xedH1szi6wKbNc/kbXxMFUk+gv
5FjmEWjAZD8DrBcqmYW3bx3mZy7W3kqyVvlnO2OTKBYyQme45hKCxEQzxH33iQMusKi7B0p8/LV+
iK250M8Lw89BvaT4PyNQLpH8NQIIUW7Q5kPGzs3qbR0dqrni9igFmHO3O+cJyPgQTyvB5puEl6Yx
1bcGYfclODEedEVdnEWarNsSTKYm1rfHTrgVFV7G0PLyhGi/90x3+X+7Sp3axedQXd9aCk+aebVT
oad0KYSDiP3ifFHtsyPx0f3ghCwx8iYF+DuN4B2XNxPkqx7KaKc07T2zSGX5zoZUfZn6s9AJigyU
QfimDFHuFccOeSyD1ZL/D/hMgIwVs6DYJZDfvXSZQ4cZok/6t3x9kbTAYYr2yn0EcsjL92N3Rb7u
ftENtGqLuRx+Uc1T2/PFmUDkIDbQwae0+6bCGzkhSX11OtA72ToXDj4HbRiMGDgHrInMEoPeen6F
wMhk/cAHp0C9bpIeOETFn36V4vMSMbdjANOaaoQUrvUXpJkIUy85Kwes8hhiX76tRpR8RIj64m5G
uKUVZAFCarNC+9TzEPi+z3CM6g4w47I4LF1WLr6I6z8PBrkZQ6OjjUcLUSTNJyWWmPFloHmaCNgw
M0S0cwBceTdAMy9gt4T+O1LJQHYdjyOiQnHcW8ds6Q+r2QAInVMG/HXlkL/5G/SqVzkm0j9+XVzm
dkw5HLzpXXFAdqjL9t/u9b2foVn8flTB8hbEgbJqq54+LMqAkFsCh6ModrwS22rF/jQ43URmacVz
Q+eoYUeFIbO2CPDpIwI0ge86D1d/W9wwaJwShngJ9QWMKnjA6KIi5dg+bIiLht1Ei+RKtwEfJDUd
PDTENLO/CwfdQUikWI4yevCYUBZReG9dXlyCdCzwb3YTdaiBHCHm9DBIuDqR2BLhwuaIV9Qi05A6
qB0urHFV8cFcd7aRasUyCbRCeD7rbl8BQ8zSE+imOzsxk4pOjqXjQE78r+MTGc8qHf49rz0WIe7a
7qR8sV3Hs5E4wox5Bi0l2DbioR721JnFAaEe4GwHMmAmiNMiC5DTLcZ0vRVgaVaoh9ro50pyKc56
iZ9DE2Q5TeqNriBTsFJbc2j43hnQ82gM5oagqLAztyQU9vLOicwOgYTxo9+sNBckuvHagx4tTJ53
leobJQG+AhT6c4LyhNaK+bYB1WBEn0quNcaHEtcjPdVD3m91OUBSRkTYarJajhNRXscAey751FhG
DPrF2bV+2FPreFkaV9USztFtzphPjK61IanEFBIPggW5a+IV5KDN9aQ+WrCoNIHEBl74nJmWG4ie
Qle1ITGzF2OewYKuaidDoEVzONmcEKevFHgi0gvuyvLo0mmYmk8AjIPozYhPAfTrrSDMk/pR3m1M
W1OecCLPdDMa1mq7M6rKdgcYAOHN/tX47mK5JmeY8wnjd+VBQWiZDQVdH1idAwr8pgEGfKGIgYwD
dN+2udgyqHXk0nW3r1PVnoJO1bUvOW0doSnhfZVFzRwVfMKeju03+LVXzb4wV1Y4so+Wlr4YARc8
DD7E8dr76BKD1FFG2spUJ2C7FZhzpK3Im6KxA1iHw6Dz/XMeJGuHaciQQbeCH0hkw12aPX+w2FLv
0gDIQZrs16My5SfWerhf+pWVuRfJTtumcPOQffvSEbzQoW2jFjp+l4FgTfUIR1o5sQ0Zxpc1MC7i
NkMcnYFSH5nMqzJwxIvlxlvaZzUsmiwQt0/Js7vJEuyRF/erUUbckKACAzUKScw4kDEWvobwqoSq
JcMS2w/ztiSheyl6/dogCD5H3bve69Djs5zsPdLVwYSPqNinpRE8Fb45VR3kjouq0a+3ZzdvLbEc
2fLfLqtT8U3GYpEjX3oK4/zP3N/dtN6EN5PW9hnyHrK2B+Hyq1kIdssreiJr+nxQ5c89JoPkHDh1
DlSs0Lmrg89ZbC7qBx88rix/kimGBLiJ0dWiMVDqIp71K88lb90EXNXABkld/lIVDQ1nxdDZm8tS
pp2nfN7LbjyrmWQ2eUWEuC7L0pfe1verPY+gG+SpB5hSt2CZ45ApApQ+URPPehNJ71/rPye4r01g
d1360uzDHW46OZsdMMHFTP3bo2o9OeexWqGZ2KIPpzaItKvFJTEe+Qmqf3DqpaAMD9pu7OIEQkh6
hG3ePFpIO/wnP2s2bFgY7lqQvmS1wjXxvhMJi2Hio4oCPu9TscsnE2lQKxfTYDnePWDP/r9EEO4P
bY9p3aRuBDHN4lTM4q8xgExcCI2mRHy2xhivFqCui3bN7bX/20hZLDcf4CaQI2PiETLFK5eotQi7
WDaD0kDdlGKlk/Z+zE8axLEsvsh3DKbKHjHzevbDPSJ4oxpdgNA8RnYkV4O7KZcf/9CMMGB8zcoF
OKgOCeaOd6oc21QZ+WqE5v1EaYE6KQm9TCVaHF2u+p+RxgJ09ALX3Y4MV3QcNbEUIcp1P9nD+cJw
8I6ZWmAlT7eH9ZYzvVpqAGHBYERsXJ0TdfH9w+9R+UVEg2jYTNoeq88j18p6IxpjLTw/AEp92lXj
VrXngzdXF/l1jVhFeBeC2D9I5F42bFcYh+vVfjHC3jmbsH9WFbwPa9RvFtC+Bryccls+MEHIDMx7
qhXafGNj/a+KP4Y+EF5jdVoO+LqcE/h84C6qHXc/7HgO5UVl8x9rI2mjkES8iNsgAGEchTuC3sTA
nW34sCD3iczCGPyfQGAUHQ1g7X0P3llnsQ5NI4KDjJQhATqTeDD9KGfs8mexUViTr+Difs/p24gX
9s4wS40d8rB5dLMif9jgEU4NBBS4QWHFtKPN+nJyR34dcnUX7PnTxPdx08SicSfmGMAdSPP6xw5P
I5/LYCe+u6z+A4qW+G0aqatfhiO6XW3NJerco64ID/ndM875l0CK/rc2aHDD7imNPJ9SANWFqIvl
SwBO19mYAdGWSZvKhMzSOd0BD+c8qNvw2gg1Iq5Ytkzl5Pkmi0qRQ9BY1cEZLDTnxfCjj/9I/+sf
PyJZqPOwPCOxllhaBrqo2O4UYuMauHdGFyO9bIZmZ/vHkAmAKKZ0IyGKRK9R3M5usIB/hAtWZCo9
9zkE5CfCv7tnGRnuNohBNKLRDjLYSKs5ulMq6Eg/P0igdvfUqgLhBAZ2DgwUQ91A1nWtXWkNEJWj
/BX9pyquDylip0TZK7FRtAhBMQe7QM5W8mrdnSib4DeH2clqOy6/c524FeqDnwq0/XZN/OBsdQzU
gDLpFZWIGiQ2QdLmtDSqSzcPBfnBMXIxAYTOMqbCVJmeurj2owmGgIo7hL8iMgN2GDdmE3MbZW7q
LpWo3lsIXJjh3KIc0WjaOtFaCtjTNDdo8VLsOLoxRA7idOBSyvo48v5ZgihPEwqofTrwOx7zSEGP
Ns1CNbXozRh0Gy1wty5I3W1zUunoHfdA6rl1K5TQROfhO/CuHmefTc2snQphjzXyN+xoG5p1MdPk
uXgLjMDGCcxC9b95DhpfjohIEMmPsMCvfYJ9Chh8bGH88iWyci81Nbr9cVgQOxssi5zWx+CiH0S8
9BjOjyE0yyhlSEVB4Mvq4l5gFIeyBNi58GEys6T6aTkjaYbOvvdrkRIT6kuZKf8ZSz8trJBpE44s
tvZeXNrb4RPNurE/Ht56PSrhA07JIwXCW2j4yP9/p/jlFpOLPR/t6jzv6ocOaIoP/xq+AtG5/WlW
k/w59+RcxRmB4WsclnZqa8CM8jGC66eUxx6hr73izX7mU1tQt2taUvonsdW0hAUJ2/zNSesBLTSz
Zr7MpRWYo3Oe3Z5xFokA0s+SL5+8ALJdqwWyHT18c6RXpTYin9XeOs2zsgNsi5h5/PW2d4JydrxW
SxvJFFEe5r4hAufIyZ2LtRu2khLNuEPoWnFL3H/6vA3tC6xfqi7CwMAYAwaodZ2wNOeFhQ9cupyW
kPQA3WlUvztJ6DkHQ2YDEIFNbx4hYwT9mVfJdQghSbCkN32tuhwHZWvbwn+cc0xqoAkaqjJDKRgd
3syz4i9ebU8s0QVYlVR7WixESTW9EzhoOoYmd6eHnWFCNoaRvBIuI23eCPClIH4KMwfB1yRTrpFO
MrdpwXEeUyAuoyshAvFBgNnkuARu23KO0M2hPsT1m66WgOTh8+TlXa6MXcoTIFXt0x8Ouw/zYPTT
XRQoRlNYgq1s8/d3a4B/9PrwIQjZysQmiDVP97hXs46YJUmQejdWrIj0ILiDxydxp4yCmqyLZBaO
OcE+IFE8z74gRCKXRuOIRXoYFRaOhRYcHUi5iN9Tef4G7cLAWoPlB+gj8yoeL7q3M2meUmZUpnqo
6vfmyDlJrldacCeeHPcHZPz5BOuLdXGFsRQEeO5IkgR3pmoDe/GxK96IZnTvoakU/t7q2KmLzbUe
ba/Sn945OOaZ5VrTnEWB0IP+8MhCCdAq0X1qIncKYWYk1wnXTZ6jl1heoQkZAh5eapHBurLIXO6F
32i3eFguB9ZoVD+d9PUN2eNTTdz3guHkTOdDMRR3lY3aOxs1BIJ2KQMmyOOkOZd0UeeLISl73E3d
Ss6guahT/JUigIp+dV/Zhio4qPTyXMVamE4CecH+GGigVxf8t594xLhfMCSmazumQw72p1GfI4EW
GIVO+NRK8jw+sdg7C+ioKv9toCqyFLOAlgoKeG/4SMNjLG8CsBUR4HA+3gnbs6xxkY+kSdKQeOlu
QWMNc3VAgpbMMbaocgvz5jFxInX2BBOR1R8Sngl+T1rrpXfOMr385acd+5F2Taa4638MX1Qb9lUm
J9SnrNJiubRhN+u9mOBx1mhJNoye2mYhrVYoXMM3DCQ24SUGMIinHNifrmoBZcQ9n4Ylh2Ee/WrK
5+7IUCFZ7FfDKTLdbsTX4sgdPMCc0vwiUuEFpAaTuUG30J6eQrFgu64XR3ZlDq+Y/j+74niZYJOB
HjxpSYikm87y3aUkOc3ZSq0wN3f1sh1bIZb/ZV1FHQyLvHqUhrtHTeLXYcqfyCL2fKYHmaPGjaBc
BnSYFNoerJ4zNFpaYg9wo9NL0RcUhN0sQq+Pw99Xmx3nBgFaENJ8Y4i5Ns4I2giWZESWNPbV814T
yshhc36tD8O519Ae9wtmsJPpTHaSe/ZVHHWz3MT/ImlHOG7fjwII4W3fjTdTnDw5e8eePFqYjg8S
TWlyclqr7263sVjCZSkKldyKAo0paPZAS20MEzc9OS7X9XOwFBLynVlyTJ38L5SqVN3Gb5tFgIng
MnLN+uSJsZLyRe9IjK/Mddg+t+C4Zejf9mX15VBPO/c03cC+Jp618uAfZJ6yvGeXJVMZNU1ywAa/
JxliYTaZhOVKUtq/bGzM+oWqxKW7NKcOlhpO6W47AJrpWfKsJ2XTaEZI1VbQXYQXDsc6y2J7Ns4I
gSZaNHXIHDx5VpLFemV0iqzpJugh87xeEg+rLEeuk06/sYsgZTzpI3RyKq8ntgOXlcOCcTVrmEMj
di7mFEn8YZSFXyt0lYSCHTvjZt/9PBaK/4+IHVF2m9J+BjVF5uXOBdlLCCRc5kH3Eq/fom5cQKnB
Dcp6IG+OUyLtVjyp3oMMs6PnoslUF4ip3Jia9+Y8GsfsqEdCjnXlCPa21r7Wa0qg8f6paWgEAw1i
E2lDuCC7XMag2bNv060g1fbMXwmBR7dvUQOOzZ5bAtyfYp+yDzOQ4lR9NreUjG3ZDWQaPEwAsmKf
ob7D8bas/11308kWwXKEEGQzQXos41hSy76Y/YhGKaHlWX2u58FVOZq/HZIqjb1J+14wdDbrrQK6
7jAZp0yCe5M/IhF9j2iPiyd+tG0jRRUXoAbryBzSuSzOBjarpG3LIDi6Cwmq58z7tgBc29i04sX4
7/2Di2/57ntxaxgLP6Gjytd94EacgTAP+zBpwzurwus+IM/6gVvxvDzaBmlaD08sqeK5vKeT2jHU
rSt+GhQahMWTIrAMsTM365quTgQx1vNyYqMWaHxUaZugiCcLhwjJkKOq4spHB6sONYUovBxkning
/uL20A+s2VUujI2ocKw8/E/g6+Jxy6JGJTaLUcTwxyhhayjHR7Bk9x8mJ4z8E8JR07Xf0UAX9D7i
Vvd+u2FEZ+2iKDRvD477jerD2KxZNF5VgAKsXZKwDvYdE4fFjks9hUbBlJHinjYH7ppWLP68GlKJ
/XR/5uRR0o6EHs0C7L1rJiQCg7Ow8ZsGvHbK+6NodrgLcLBzb6JS6fCAzw6FPW4q8xyFxrTgwDCD
ZbPp0ZNQGHhoNyUAroLQNpVwQ4P8zGSWY0OneSxNSEC7KVDbW195Gp0MlcpmtyWLSJbndpAlZH5n
8TWuxurN07m5pPwLu65VDMtTNLLBad6U7cEWaT/TupVzMP/QOGaKo8SPNkPagG2jNGekDXqsIgbL
Af+RGuUfQNSRb7zdgl/g89yhCkZeazJs4xmxCcf7QCzimNb6lSCPoRwGdaeHfVLGnn38yJXLnTea
WhITzHLjHq+XZuFSlGDV+j/5TefJqlywOzgvRVwKFrTHpfO1kbCyK0/pMy32UNWuIQ4w38w6SuiJ
KcMy8n1imoaFJUsFgyqoPXzIfHI3Vu1hSZgdCu1OHhFbEocpt8Lo6KVfQyzB8y0hA4RrHW6xIaQy
MjkVkh/vVcAE8zEPbtszBNFNYv4aFaQY8+mSBuTI2HYWI67nsS306JAiEibvH7BjsCRcy87zcAb1
dF0b/Dm58NJMt+DsU4c7EpW8gdGZeug+3MU2dGtUT5aIK31Tqtws7jUMAMriNmxB+909f78bG+P/
ETVMEX/X/2U0+2uXBlkXjitAVGLhhbZ+aRqSvu1CPUraTNzOzt24ru8DCZji2whukJRFk3XLogxb
tcpRmTsuVwVu9SGYRf6sBljElY8Fq4SlRh4RMgrl7JNFMalGWpZRwrO6OOjZDXD4qA4vhwhQUk5B
2ECU77iHwlNr2rUrXwBhBcWkK1u4etm8yKNRzb2CzaFRGsg300Ejc6mS2mYKavScq6GHY8iCJi6h
rF0Pp5RJFWX02VEq2fkygAwzYbgI5hVlYNa8PWYUP7qzWm5HN+N7hqQDARCUXd1lyIq7JVxTF0tl
AU2hWvMooXBOjHhNO4YNkUZ2lZChLglFn4ZUFz9ycrP6w1qN//YO1SLSNyBrP0tC44sWHDXjJj9I
pSe1wppChCaMPB4+USgXlgOUyGkSocG7ddXJFsHOo64/ZDPUP3obOndtE5oHNxL6JdqhexuLGSfC
/CidKTjImWh3sOVaNdzyqRfPerVdziLlE9ROtDVHkZNmIPFjY3KCYfXphSp9avz0cu8LzlzJzlGM
hLs1oblyRr0VpPSO5CsJOOPJ2Rv5GE9KP8+jEqkyRXEjLWse6pkdspP7HuN3Lvwj3KIScQDQYTcd
xl6GEUSU5Wfepla7JSlIhKgLbIX2KUbvlQpXhNVVoUlVab8dQtvxv6tyvVhgoaqLANVnAJINvA6n
krcpaSGlKlKnl69b5HXVCuHlKGZ65hizhbWxBuHydfnx+GPmXDLoFeWnH/VyeIr59Y2VH8a/uqpR
Zs893Rhw57bneujsQTns/n0bqVyf3x459aodF4JeR2tpGenpbXmd0wvudIvCE9eiH6E8K7KTCPpL
wKAbor/PYKHOKVV53+/yntm0aPdvsc1pATWT2bzZr3QcEmWtgvUuvGbU65zl1uL5L2GBtaoYsxDI
v9MXbHxqUiahT6TNff8X/3tFONDfqGLj1f0qgqWgQtqmTh+7MFQgZZRjfdbzD1HFVWWDEbkgX/YA
33O+ORcYxhBo4KkxkZgjwI/WmLEDOdhOb/cspQ4SdfjkF2qL5DoGwxl/eWCXRiWqomaRaQhsAuoj
6cckMpnkvX+Wsb5di8OYzs45TH7ZbnCm7ksXY8BJvEiOsi5VCKEN/rYS+DfOdkyrOW61sEm+4vng
eMxk9OZlEg3YBELj7Zl0aLU7Eu51XRkj9D8v+Lm1uKSXzMk3H1hw/oe3RLuaQ6mqEh79tMUeypaP
gPC0/l8GRbAfzwrsGNG8S5fg1dXizLMDf+I1c26/SAYFmqBb9Ax6hUAWEBHBUy457CCNQ/c+VeyF
atH1s51464gkZHUz8sM9UaujxewvCHnfLE++RTNz7vsQJ6knMvDWExQUIPO+hRQnKSLhEYmoeDJ3
QvC6sZkRfcGgi32cKOxhc6GNUiZQ7Gw8ZGR0dFIsl7Kx95x7F6tAz2SD+2DOdJoN72/fbbtxqQ7p
VzHt8RqDNVewcIV2W63PpB/zGfVKHDdkcc2GmcVvn9cN3qkF4EREvJVl9GDZT/cjKKuK31GWR5oc
mHvxLThvzLfSBoeG6+aO6HmqqpRrngrpXTn0VcVRbA3/llVVgUGmRLRXGm4soBFSw0Qj91Cn52mn
TwTUYUKCwqCBAVo0sNmgANtOVSLO0a7ICXTuR4Fmvu724Km09dMQ2Ii0kGMnoEd3H6s/Lgj7gAU9
CnaHssE2vRsBaWIqV9EKDvers9iagepNcDJ/vSlkYcabiNwZuZpcEbAhdj0CZgkFVfL6NYO2vjAA
LdFJ1KrhRCsHCmHgeZiTYR5qp4FVynDia5WkA3xObsQW85KjTWd35/It0vXlPZAJLul9JP5kuSqY
vmc//ByUMqBoBBiPSmYh6wsHijcyEvcp/ezNxFYSSiUsfjDMTBi2kqozPjSrt60n0XcRTjWWT9a5
P8rOuTjyaIrg1eyIzNs19UDWpc3orYBK5CgvcAY+BDBrA1PbGYdU3sgYpQUohj+3SBvOo1BWRThU
KKaL7E3Ayp38w5w68BUerNhFNAscx/5aXCj1vkKM/3/G7yDzYDBPTjRUlTA5+GTZ81rfph/UQXRA
nMcdA8olHj7XFOMtIwS4SVSKARASs6xOks0morbc1ImlmLoLevWJP3WqM4Bn5XHmrYTjdCkvedEz
O+hNFsifzrhJPrFSIFR1UD2dJYGcuWkzLBSJvzoLeiO95X+/8inouQoNdYHNzyjQGqFPDjSGvvoe
eMvfoRSqIhsI0a5pyeP7pzvz++K0M1wHd4vQWRXfGeYttbTF3OEtZxmcX1iZepPZS5EvuEl95ydk
SjJH9ClRJfBgzepmqIDhGjQssw+vaEuU1SuhBMMBgu8El+OKvY8fmyAXnnF3aKVPNePw8kg8cDvP
+ZphcyRyhxYPU88PFKG6pMjU6dyAkPx81ZTDlB2EPKtYYAO3Q2CXW0KYNmXWxGIH7vaJS7A04M9+
u5ZIB/+vZZPm7ss77NOEI6MZMMTnH8wNc0BNp/oegF8GjxTVfcOCWRFsjKH6TjZSokgJjVR6z4eQ
wL/d4DK5nFbOCogq/3A41IFMEKIXuXeEnbUNb2/4sNIif+EmFeJSbDJijwDXZd31ZVSM/RGr2IeC
Y4oMaQxSYgYvRNrLwX8/dPmh0bMIwmfCzy/linHEovQD0DLzy+yZpLRicCW03i7vqcpyCYCnH3PG
QsPx7WsoyJNwLiv9QOXDp308RRJXJ6tiOel+0XmInKAMwSHXfBSMlwaS+JFCiDKVQ9D/YY+fJOOe
PW2tV/60Dx0EXckdhmuAApXRNBEq5DHkECYVY+iE1HM5P855ID/hLuqfkaOfbcHduUdev77SYe8s
/wRBSsicvSzISpFIa4FIeZN9Dc5IQ5NtOWyOfANlTPkuunchuKJFWjd6A3qIxXdYP40YEyIf9c0B
4APUnMPwfiH6IG/v8Bwj0mvXXuSNI1A9ihm0B+h54YONflC+5CsPXhk9KQFW83eO+55aVdSQlyJu
Es6JSywed8CEnztIKpTt2u6M8Vf7e2b3wQZZ47eu+hIp21bbsuR9IJwrIAbWHCeO43cTAI7uMb05
lbMtCvO1fcW290iodvMCNYexvQkNbn9EpBk4a2kyT2dbMjvR2Telzhp/drdYq4A0oTyYvzn75NT4
RaWj9pVjidkcvR+ITuei27tSUAPoU7sztY370hCNoYnNKRN5WO0bAxgTdjlnZZBCMtoUMmSq00xI
EuTp4oi2Z30QwsU2rWOC5UA+1+BvOWOe4IjXUVBuPMg614/zitSmh8+VhwSpc8roUv0Map5TWxjK
cLIzoDwLYCJg7eCoVN7mcWUgl3gr9SlfDtifUELofVvup/nExfmwrSSZ+sgxhAnxXW2j3CfcIm7S
kVrN82mXPN6ZEEhrTsBxBGD16HWbN9kpNaQbrUB5+3rq4yCMwXLokYrPWLolKzVTq3tv1yzqzFkb
pfohbNle1/paPKGKtcXazWijVTNHwpeIdgIhOO2snhIq3aEJB3nP5XuyMDcO5yJ/HvlX2jvUZDFa
TL0aft0M1HDW64BHw0XrubWUdTFnAkp8U/UeP72u5W7zV8lL+m5g0gWAa+jOSxw5hHlyfCq7cUS/
+VbDtrESEpna/mmNtMF2ekuTRxgqK0mM5+aS78qOM0rSMvrX5jyfGcin1JMLeKo7QTP4v+wpGUtK
KA08Jz+kF2/FC54t0Aiv6Gge9zfre+AvDSUWunZ7XjPcjXgyL3Yj0o5pR4JdqMd3yb8A8Ed6DRv0
Nzth8hb1JFJTgYMUVfnEX+S45idmtS+2Zl55b84giNiKbsPXgLogvC8lfT2NiR4iWVFNtg0VpV3+
lvuEt8A+/SBSJvJVbVs6rkhkDaCOErIUo5ZatQB5xg2U++dK/5n1szr0fMaD+EsMqqAAmSK9ul7+
dSnyyyhTNl027HOkPkE4WDVh2D/mURtYuhLildAX19jw1aLWnDr2/8k1BktNrSqSbZtvSH5UsX6c
ixJaTgT3pO2WGNUPGI3KsTLeHyst3NMTIh/HBGNYnKqwwt2G+435bBy/sSjhq2ycXmbegR68ZNPs
NKm2RUQSzln7ar76eTI7EYicMzJzJs4l4XQrrIT9evqoN9etw7Y0Pwi9hLCDBNhhQ48WfeIwd+F2
HJ6/ezuNYj6skXdJ6mQw1IKHV6+wo9QZmZsKDWHonsiuzu4XZNvdy+Gq2549khy+szbCuitrKitG
9V84Lc+U3OOcKCrJSJQ+l7544GdgGzRsHTWSgKlqavrLccVznG2X4/XLR3H9p2/ek7ajExfaywdz
eY1GERH/AgW16c1Bmv9wf7i6jDuY83LQFgvRQmiuVgznGBFKmE1EJ+tz/s1Ea/NZDLlNEX9MPpCp
bCTSa3VZ2KKTS8E7i/+jJrlhZrjcA4pcHuLVvMOsLK4gSZvyKJQsbMeEguQXYY50XmPzSMtAP+Ct
enEFT9diRMF3clk6APfyVXSaB/MS9kBYe4rq3NoxGh0hT90FbGwgeTn3klo/SWsVVJ5/U3xlDgG2
2ReTODcfye++B4GOyajlvwDgItqNOlzaPH3ie8EdS2W8JRSu3yc0FEJkkFkv6Tdhf6Hduxljf1Vd
w9lnnXqwuKeaf8yKTvaiY55QgSXLeABWVPodPzL3lE2JEC7PbGRpHdc95JvUZ29wAJ6O5Jw3UXYs
YMjDf2F5w2xo2UWQnT5iOJioLrunTZBOEL8Z+OsRVewls1R+DdcxSjJNpNJQ5o9JXxl5AO/Jz464
siTs1eWJlILuNZr2afGce1l7/IC5HEWfvMVVCkGX0OrS/C5hUGRX4skG6EWIeX7nUK5KbiOHWx+D
waT4loxxQ+5FCH8LgeP520SWNN+g4nffYbyR/OVDSLAan86WSrupAvE3FWrMvFxjKLKcHNjsk3A+
27mdU8DODYCVRojMaJ3DI3wH6MGsNISrIvE2ZmD2RwGHF7egkTHXYPfvRfyoGbVbjUla48wImzg7
0/bWYmVAkgzSLohdTLE/3C8vSahHcZUzVFTeIGXbC8sa9lWMO/bDrpD247MpY38Xye5d1a4MZfLj
PXyqrxkadwYRyFeoLMIeb83MM3aOHtI09KR4UJ3hyq2d9bJVP8ic11/7EhFecNxhjzkYMenmH74B
TFSEsBvwk8317GeVHc/hbMJ/XrCPfdnkJW3cYQZdK05drYqwtmXczUNXRy4EwSdoBkxRXdh039oj
BvuQaWt+fYq1TSZvWp/8kx3S7kKgdLEQJ41GvscfBO07cIwpgvGXWy6hXJ4xQmcHqkRCs4dIZJiy
bg2iKRWW/jgQgM9kOBc2NZXqCj9Va7eycFMFVVz1vnIOpTqmau9XZLozccbk16lN8ZuLIBuMvdGz
Z7LktsCzK5xa42WT0YW2Fk5vCCAfzHw34yIcom3muOZXLXRjZ8FFb1a21z2LQOTOJYynVtg9pR/9
4oUFU0bWtOpaORB73M8eFjulxeApKhgc8Hx13aNXJQIXAClz0pjJ5hvvPm6eYXnLdlpZTBr8jC1I
6kAiJpad56TwvHcNC3w0yDctdqLjTDKxkGFiikwvv2bEsus2ttNJfN2Z8zTNbXZMkp8z6j8S+hYI
EOT89qvtBW63KNvcWpLIOvVYW3JalGGXL8ZzhHn6bKNhnouxlYLJ24FWLFS4fS+cczsMkkiBfPoP
zMGslL0mzQBPpwXaHuKw4SQJ3jBg8odFZdtHOzEjyqLlkSMXmxv6f2hqZeTayQ8GMyGrWhnFF+8P
+RGr9gMZuDupJ8OPNuyM/oF2E2nnXfeJ19FPbSBT+7esLAhC8O6guRIdzxjIS1Pwn6B7X+GLWc9U
Hlp7ceR0uwIe6AI76SBJakuiyawRMRlHr9RAGv5F5QmQknJYPITW9tThPickPsYoy1pvT3Qq9Hu5
+5pngthwaSZaTa0gNjffiYCHc/QcQfSQIuUEstiGivaI8FDrd+rH8t2TsKLlYGIHeRnlzhdBhH3t
fbQ6kN2JnkVJNvy82Hiby1/bbcegFNjRElkSesX8dIB1oGJAXlMKVE3FLudsZtVqEZvlzG1viqC2
/u2ffBG0FmiNb1eKz7PFlgPwgGqwKCO7NrI4scsLxIwBKGsM1eafWcip84A81G8wdmnfozJRpM1J
kfpaRH88tzEvP7Ho7pHP1OWVwYOdVhDqaCc7KZdV7ojU0VzVxeM1SKQ3apOlHolXc+eR+E4lV4ep
NbXp/JrmTRqhf1ieU0NekHwyE39LKNSAwruMmkLFCvqq2dDJKFDOymBRKr7AMmJ2FREby84JvY8K
GHeD/aZDUv/zFoGpf1RJ1awMzDdJfHWajHknig7QVtC3/qu53QDDSeswTO9K6dZBV0idqYH1HnXN
DngHAz5oy0RxOIHxFTGf37In58U1OWu7WmM1lMCeDRnf/s9tZ5QgrcHRLj0NyCG4KM1852uK5zPa
+i86Aa8+4SkPchvuAopFwcY2tltZxgbLK0VS7ym6Ko5YQ7IhxTnohUkkDnP4sdrwwOqHyPu2P3nv
0ITz4ZDlBEFTjKsj9amtMdqdbrf457I/TAnZotOpwFJZRKotqilzzB1RhLTAkvzK5sfnyXwrijTp
VtRltH+Ki/2Yc4YjXV3tu3MYpDp+2eJQyzB+Vuo/adQYm6w1jN/F2T43wYCE8bb4LdvcEOlzAKnY
+kiMqTBi7iYg9yFq6iAmPf2xl4tfJxpcYjGgxjIjCoUvOdc4V677UR5Od/qtT2XNVZaLX5A1IP7j
RcGihR8He1CSs3SVkOC+UpPa27F+D2fBZjp6WtGF29tJrlrVmEU0F11fttD1HS2Ybr9bqIg3O83j
bmiZ+lamppGps6XxdsL5B0SfpVgho6usqF+G+hCCyDsxuFM+gHD0cxI6xBhZ0BxEs56WTzgkeZSx
oYYYZZ4RcwAJpKWZO9SKVVBn08aohgRUJxvpxuAZNMRB0QFhIXTHegX4/vmzHEXlBtTYWW+xV+RN
9S/yrWsA/d2W8bq5wByzlBkH5dzQuIi3W9dODElEwpI8gioIM/+ekQACM0nDOYfzXwgjSu178AK9
LmZckIrzrey+X8lA2rFSYpIkR37ErRAqECIXHcGxdLcmHPMvX8AvNJBqAdSyXTkzJQBp8GBX744n
53Fw3qXa6bQa2iH/3MYCkEV1M9LiowQLNwFZvVB1ZewWl+u4NgiS7AoxMP8QqU2BGiiastodtwjp
as0Iieshj9kaQT37WUzdsFql78A39PIJH02GOHy6wy7hPFVj051e0DhSkExWg8qI1ef6RmfS81bW
zs9UwqXqw4Z6XGV0iFGNyoqZBGmuoxbfbg2U3sHvxm478ZkfhX1+Q63sNMcJg9orlYtSLKsTkRnt
Dym+JcKSCnuJwczidNX/WwguGEhwMZHxrVouHZt8zSvjtrxZDoNrH5jX7RO2fBsuFm2uVZ8K+RrZ
KcHzBpvT9ZD6Q14JINRYWIHxMg0S//ZlR3rQ2te6lFQGPbQ84PiYmrrgH4C6V5vzoTeC3aYUr7F6
KqR1b+iE0PxcfiModLbJpKRu0atjitIypdspn39GMbKcGIcw7auQSK60AaEmXbwjsiGIYIXaxu6M
tGsrTN9uvgrIUK54QlaKw+LIojXpCypxgDOxb9qXFf0PhfspDVo7i8muaXL+JL+TQnDF3LxEzrGa
9FYAGxp7bR81mrMFDamYO45nOyqK9xB0A8tmM/947eqlpaY5mcdwf2ozva5ZsvfQ5dGPSL8cIEF6
xtNRYD29kXTAR24wys/hwQHow6IpLSLXoalqzbPfxozFzUOfpp8WFtftMgoOuOrcj5E8+Msli/CN
fgxC7IKO/OOLU0NH0d2MAUtsTS9STU3c0c1IeC7v+pC96u70E2jBSGJw4NHhKN7FLbVoWBDQaBG/
fwPUhvKd+9IPHh5bZoO2sydOFUKtIzVQkpA2GfDDnjuwEH4F61SXYgT7thePf5liVLz0iQfgH6Dr
shGRPWLDJANGmfsnXFEl9Y/O+wt2wpBqZq7f1nmPuqBtVTdXS62IaMRT8S68GgjfK8muc4GNFLGI
83KVgHyclyQx+TalCvl/VoAv0906amUqiEavtHFQBxC9fY4kjFlWqtLwZOa8DfTg62wSgMeYsZ4y
wO64jSSFC76vR9HaXw5NFiGeZVag0MXY1U6Gdni8OhgKr7Sd2N81NUVbBAZMyhPQgA01btQctdSn
LOnF/YkmBWXx1QU4csj9c9pc46kd9HzFynJd/4JEpzxtpCDv0Z6iHG548XuRywI0Fv94WPpe5gr6
T8w0gkpVQ3tx+jbfGuQHmeNl8fx0P4pDsftKOnPmWJnVDJWqIdGRSRvvae8yB+GuUghLIIIrqL64
8cJ9/yBnFQpU1IJw5iMQe+69umQNQKnCrBH/j/3hwz9biaxEoE3OHYdd57wgHKLdVuawb4BZtpfA
6kO2pfUC4+wqJA9xle1h8ntdd8CZtL0PGHJ8KnfGNFuXoZGB/C/d1H7EpxCLDlQdGbcoqtzur5VZ
ugCMyMLVNLHrxnxxYiv/a3+NxoXdM3plwXII/3FCckLlkH7VO8HckW72gxCeD71rmffD1sf2ryfu
9++KH2vPaLoBuZrBR+tYkqbkXYapGN/8c4cn7uYmLX5Qyfh+WZbZxjLA54/+G0USYp40lKWZYsjM
2tV4rbv2OW5CSkGwgP3eLUoMPPHKk5jLrcMZ/Nsmhxm8faYjwPTul80DQZWMswgK9TzysLOrgwRf
q4yWpNd6bLEHVqVnaNsT3pSRz2capVZ3VSdqe2sxDEdl7im88iEgTl0uLrHuPc4huD55hvKxNn45
GLC24BdRhK56big0OhJbkFNbJNh7Y0qvtcKcDAFCDq/eAP3kyYLSU2GjgPNez4239F0vtNyRNPpc
8AD0EFFZOVpGzpPHmRAo6CWykLhsRinGI8SX4u/HX9xuO2EwStkSIW3OMtT+Hu0PD6KO9GSNTuPL
nCvgZaPoWDG54OMaINrwQZ3g3vy+eIvnpmfJWh+CPDGJIeRLOB7TFM7YOhgY9/C2p21zB20t5hUI
sW3RlFg0yqtG26EO7J1b239Dcn4EhalF4LjzxyGn8ztLwtvdpqECIbPuW9fCmosYwbY9ZYB9cfw1
plXW34rJJV2ENeko4U5KYcw5rhOKyQG+qia6yxB6E8KcclzQFnQ3C916oWA+62aEeaM/KVt7alob
9X5VIt9M2r8VlQdJg2GEvLF7mqCGmVmXavNiHJ3z6XHprUYs7/HqvB6YJtBXyeCNgMYYroPAt5BO
wO5xIcuC121LgwsSIfoCA58f04tVD6zdLmAiuatQou4E5r8D+VP12FAQESjqkweJwUVZEA8zgkV+
vY/vR9s+AeqwCzpL1uI7hJE4L6ipV6mDl5rl6hokzvt0yet7qsrYGA2uPbDu3FkZSAuqrKwkSxRv
JRI1Xwtgqy5Wa3KfYNDSTLtMCLi8Ea3poy8mJ59MFvBO0QWlGiJ4JPLSgiIJ+YZDqMZ63pnlwaB7
Bg/MqoBY6G2PdpGan3DFFrv7fdT243uF84gYLVdjK/ya29TFY34a4g4atjvZfZRoJQN15jU3MheL
Z+D1ranmclkKWJZTI9dNFKogaS26ecpSPyIXC6FsIoe73PmY+1BF20st3Hq/0QSmW2eqtTU5xpzd
kXFBE3f8YMefdyQMW3owjzKTcR+pQzze6wxiNdsldZAaxmwn2VI/3HQ9vbOlC9q0Q5CacOHQYjV1
8gdqDQNXUMkQvKURn74MZqAi7tcKRK+fl14x/W217cPHJkBX0z0T8Z2cpr9X30+VhVG+Og0LHNkR
zWsNmFlkQlqG3DiLU59bE5/+D6IP+KLNchjws3Wktfi/cWdUaKZXlEeu4fDlwqbri3UJtINkvyzR
4KuWMLYyhLV6f9EUPHQCIzqy+/ngMuUHZM4d/lXHISLXS7nbsRzMFcuZ+BWGKqbkpdq56F3CarPV
zitpnDwZefqcMNzOEF9/fl6Rtu4rSphbCDk1p/p+RIojXlOZUvMjaAMvgzU7aFYPcslAskOvwLQK
ewJzc4JBv9gmF0v5nzXkTrEK9ZsWfkUEGXzOS+Hjqr6ljyQqa32hsYMPSx83taZgBsffa7augLbF
K7KSLQmsIEFvvxrVhs/ziPkz92IxCAFusrqN58wEYIq2Zn9Ddg1IKrTZMUQrb7km9ty4Kq1wXJIx
qkZ52wKGsVe23/NFYcFCIF+nfaCL1lD3bSd0ietsuT+rSno0HdPnR56So4bJIesAHTMCSYVxIV4r
cFBf9BU1TH/OjCxXnnMqk0AqzjD4SugyCMwYXMZAaU7oW/N9uT8q4pRBwP8m2hOmDgXJDYsv74HC
1nrpNIJpR2nzGs/Y4idvrLUwCqTVPYs/JME1MkZ2DC7rppIm2AgxPhM3Xip8BPg4TzCBgYg/q+r6
Uy3W5bt9jSiIEdJ7iMAuZh1ufYABsFGUUmXJ6gciqzJ+aDhe/EumFsCAwgRnqDRjtM4fZgzWEqx8
Uju4NxiBsCQd4Q7oZR6KxGwd0e8yFqv394g4yytOvM525IZtmnZL8EzwndRVr7K25rYHKIolkLgd
CnALhrgCfdbslj4SNH8I20MGaoMxYsviY3H4a7h7jnmUM8q1zngYOkHJJaPG24ru9tQ3Qhzt6gvD
f2CswHaywv3KRglGbnYQCVk8w9n+xLLL/6R1FCh84Kk2B3dvEQvcNtBZ1cDMvzzlqKlUCgD/WJZj
wAoqqlJtenlE7+SuaPXYTxTjO70eOFX6lXwOAhnj7+eCLSHbFeF+aae5DpgRcSf6tUXGlUMfX+tm
iSZepHtzzioy0UpZZMA/swrPrYlh/Bmw493xFHVyJLpjw0T2DorhETx44+qoY7CaV/B1PO2glRFE
DP8pBs2pZmBt8rg9uwT36VU/1wak+Ba3Umq+4eamqHGcpTTjHd5cwZXAspedxSTh2WJn06tS3hmd
g1r8kODSvkGgP3mDzf757r2FCz/2n9a8PlBsg0Q6YryT/gbk2UZAyxLSAzwad+fGlTVcvt80BOKa
XpxydiajB8k9v11WiVM5LLHRkER11KL1aC6AcqehFqre5fJXiwiMJO02s8EMAq5Ql/+VhI/G8M57
LbjqKdqwKLnhJca6Xnxm4Ick5M6HLNa0wLuIOqTSUKP/v4KN7xTQmVQXVqlIGkRTpUMEl949Sm68
eSjZK+MDhKTuWKFAordb6IHdLn45JB5QUWYCartR4FJ4Vf2KuclpP1FLhQWkxvFzMbZWQCdVwsIa
lC62/YPYCxGN5oBkygqnL/Ixit8ymmvRHPuxb/64PL/f0tbLfsvJSHcq36pavNOeIKP+Mmz56jG9
XUwDMrZplXgMHfUsbVIOK/jvRAJLfBl3G+TN00nt1emNQAAxeRAzDwRDpdmJZaOhhAaxgbU/08PX
XNCT6FLXxOBKKIy1w9hy/Szw9Fwn7aYP92O6dV7nOUlhvkTbZqgTlqmxM8ZprcsXbBlCuTUZtJ6D
CKm4j6p9d2F4P4AbTGCfobCFXkG1NEvimmwT7/JA2Z1r0+nU8gfzi52x8zj7aBf2li3zD6HCarGl
QGeopKse0Dri/+P8YNaooWAM+NBpOvvAQmblgDGneCCVUNe7pxxT1TDdAxIH1QVikw70uqbljqLQ
FkQ5x6oRt1Wm7H3D8LkuRZMgvT/xWqw/tFud5H4NneXr6aTDBdFQJQjczis/Ix9NHZQxcLo62wdi
Rk7PPV4iL6MAzjm858Jd0zXbLHmpOaNa1fRRMF4v0URyv8C4pz1J38vSvd6M/MOdxnMt5zfo3jgG
d3G7Y++g1cwnf+eQQY7WYMzceDyz+u2fPu829f8pVi5uKWn9I7ENeFV7EgS9MAcW8k+0yGEm1g+0
uHmDCwcvsVm7H8X9r2SSEysrYGqWZrJT/4TqPHmKgfO7BWajAOHcU4A5FS29wYJsE5nXCXU6Jhp4
5udx4rzstQtsXZrBW4fFUHmXX/1avxzU7OcnVQHXE9JjCqvZub/HnLsxCFOfMsK3E2oe8QVJhdnC
dUB/o85HPBZ+RAP6FgB3hX3paQ0fx8uenP+9CFdNcScg5bR7v3pt+1CwD0iXF5/af/cZkfLrDtyQ
+I2K3ehgOZ4/gf95nOKsZEJan/H30Rdv6m+WNjBVLYOxhTH7nsG7tl4W4onO7D5Ea0gcNOo2RAtT
pwOMCosw91N6dqRe9cWt8X381k+r+yq3hMYfk96qXDmDBzWZVdEnliuFKvYwqr6SE7E7u6RsGMz2
9++aEPWZzC+TaN7hVdasQG/ADqdd38OH1Xn/NcFEE9rmFzTcG/Fjkx2KvCfoyMeloPZmlwGwqZGd
C/dVDNwNMJH5QiAw/Q4wW8s2JshulX1KbqFjvCWpb60uDLUfGbxHshwelO+6BozubHSQC04z5MNG
JDZevrRq7dZNnmgN9miyVTUdOFMxFGrD5U0MHOo47Mi8WoJCY2OUSssqe7N/1ulmNELGwxWy/S5x
wki1lwGjDyjVVkYxWyEdODB25q6gD4nRw+r1gUkdRPGAGCeZFK9eOpIA5DR6yYTdWFJdLMcqfWop
DTgHEEQIx5s6UfD5XOYbDmk/qeA6+oa32oPF3mbzs3KHoXuam3725HI7xw3H02p22v3uJJvWblwY
1l0RDHJCvFpR7SHHCysJupaK2eEIG7EDUN4x35OezJcqsnwKg0ymVVH0rOnJn5q51sx80+SH8Zk2
QbSP3xvVTDIYQvyziis2WE3vWI1SHoLhhAR2HiVGCTPbKCZ0BjNKSeE0t4+opO9G4tW/7WjW14i9
m+4nAWq5KgOT7RxNc5CpxW8c9w2x6qka5MpaLgI9Ab+HyxUoQ7CogZbcc2YcoVPqwGlqRVYhVp5V
kHFNF/gZeaXedURSyDtyPQWO7hKc2AHjUCsq3i3Un+/pND7j7ngXIkkGGL0gC0TU9gkszMBtsG4p
Xvkd5AdK5yKwzc7l0ubNZNQD+QGLpHdj9eWwZ1YjdoNPlFLxsP4HEhYaWNMcDcFmaCVW+ssRy8DE
HXD6kE9VYfGrcwrCsYtyX/THSwPhnJNHxmNE5nSxNAkZoM9nd03fDXj/cFwkoqfJtRTqqHdK5Ss4
/MaZMHPxg9NnG8ql/0oH7oDO4JRv5L4a73OxPAr23FCwcMRdrZvpHLntZ6VM5PtWzlTWEzKftQDf
/1md+DdwCaQG/MF2ocNhp4eUmqzjhByDbVEiy237Yf64jM4UAxwxadido58jesu3GUYmb7Dclkpc
uh25VcvvA2aiERxYKq/eAt0eFTHbY1Dp29jmG4As/UmZpeqS5pQTg/LtSsIDGokkqEoTvfmSuRhU
SYaVxUyEVjKsxK9xnb6ECtqCbpbIlzCPdyShu7dtITdHbqjnxXQPJeuKewVxqdXkMhy0UbDK6a0g
TLTRVDJkM8xJLjfAFJvMst+YlF7R08qnIh+P5vhZsEAa7MvAF3I5AKTbWFw9ze0rLUXILpqYOmn+
M9l3DjBh/jOI0FRX0B55aPwF2smktW5SKDkDXK62dCKL2+ClRcnDzLyox2M27JmEso5zwYsZcwcv
mjv+rADRb6cyjtDNPeRfL0Qh14f+gE6M3XiNfcwYFzVJfD2kJTwS1SadXd/Y7MilD5oi3Ec3kRyt
iHOpcK9uHUJ1m2LQbP9WaPVkuHdKCwAWAy/1/FP1gzrVEPFUAbbrTgxm8Z+WsX9XEn3/JztAJmTk
63yPBKixL4nR0v51lKPqITlWMb9+tDTXZrav3tIo4rb1Ac6tX5a7PoyWA5DXTP16wZHlT19aR+Pk
6zC24Y5ybfOffBLl8WDz2DJV+5Q21/eK4tfomzRM4HHt3sFC8XncU0Aq7GE9c9XrRbrSQr2qhEhK
MTHjJWU5XFWIQpgbenK1k/1lHKqitlAXjqNUWohImYfl7xn2FdkJbACxSbOSTzPrnlLqLVKYTaHZ
1Gzzk1d+EOoYnJGqyQuz4IZp2dyToSWQYVJ9nje/fjIBc03ueBOiw89AfYtSN4Op3aTG4ybjKEeI
n0f/oUz+5W+c8NQMyMlljJiIi2RnSAH90D+xnnEm93TSXvs1VkRGLWy4J4GopBgHbJdq1/qsghmZ
JoiQLs3ggI0G4W3hY1P/dkd+7yYtXM2OIXLXj++/FO7CQuLsvQqn21QboPd1hqx6qwJ5uUnAEB/9
KF2si66/dYhWw5MNUwMgSTBB8T/T7haoGsVXYyA4XkVJaT8sDUa3vrlFWIjLda2Xq/wbCTC+UCAk
mElmwfnaaxBcS06p86ENyhwMAoLma3499UZYelzkhC8PxOVGSdfVoTcan6e32G0Yfk7R4tg+E4wj
3ezepcOyyN1z9vz0mf4iHUXZuuuNVs089BKIFvbRi4Aak+1fyMWNg3ZnubVpvYKcQbpDri2vrG1w
zofkRBcFhJo+TI9P0OJFGCkhOx7EBYeyrNU8dd0iz9SHG084YQ1QM2arIOF/XyUn9M2rTEGMF2Bt
8sqQb+ZrMdtPKRO1WBHDxXp+yH1yRcEzZq5z5jo54EkAdA2IpAgem8H29271HPPu4PjdlXIO/B11
gpAYhqYm3rMPm2sN7puI7VZ9hgo6W6tShqs6Fq7Yi6+O/j23fSmIDB5T5tnvLoWiw+Lpv7fdUXT8
+2ysq6lKqawCO1cM2v0+y+3ZXrcf6yXUCa6RSUAGgx2HD6JkcsMIWcBOztdBBBR+ka0Nx09MYL2Z
ENQHmJ+OxCU2Z+4Adp52WzXNxKwPZ2WCsLhLXjtpeqAQBPhYRRYZmQAFWK3+3yssHWZcyKSUk4CH
qZLgeAbsJqqqQhy3A/uaMiAqTbOGoK4O6yBHnKEE13zGv1cyXOjOrBBqfxaqS2DxIR9PX2qNt4OC
LbZ/JLpLi5MUpvXZ/5s4W/r15QRvzcozfBOhpKo7vYq+mGD0wlfUKjM99W08ivxMzwOSxuehfPwd
N3TjvmmMlH9AOCbEQ8+uhc5ZJTbahBpy4JVxXoc66wuSlWOHSsXoo8ldk+diPtcn9GKYydZTDPaR
A0SC0zA96gpNR5RF/F7RLLuCUruncMe4XXmRqeIbWVCQjwnjcIIoP14G09xD6qcc7ZDkqYlrb9Rf
NpdgLBxxNfFLVqbhgy46+BLlI6LEgAVXDXEH0CZDZH2TBanZvXAkpT/x8YEYFJxhrOIlmDIUAR9k
Rkw73ATmF1QsoEmT4mDlCW8BY437d+qFCYhZ+rMSMOLetu6gnOu6TD2I5u1LXM7HVFxyHdB8xBMC
ogDl4cfC8ghwa8iH/Qolc380mzAsGwsET3oEX3/5aK7Tux7YOLjup08y9QXqxvjTuUS1NW0f0iE8
c91M46e+tYbigjE4oYGYfVb/6Gph1HdbesqNnJqMTCLlKvsZdZrtcfOFQZ7UNAAzl8oZkdiWv2Zc
THALDzs8EIhmlfKWDd0JU35qgEbNErCG5bRY5TllNAr02dWxOwSHVF7dQE0yQyOuyObV+s7nq09s
m9d2uqKiHo2alP7bNSy0LCYZqqAJ9spLU2QLVbQOrUnky0ZyX/fpyK68MsghCz2zzZulNghq8v6q
PJb1Tm22duH3UDOe92pM3HBsjoB4KPUS13RmHA0pQWzlXfGFZ/9Xqc7otMD83U5hnTg++GOougpr
js8U1+O6i2ZOv9eQggl2Jz37L/xGMop1lgAJs2x+YUogAyQn7xBOQ2zl7uH4871U/Gcr7FBlMLfo
udpoipkrZCfV4TkUaL5g0M7dateVSRvHQ1Kwl9EVnj5ZMB3t3umzy6qmnh6wgvrWuRsB4Y792k68
OjEwKOXMhrUakq7Je/SpBhBMnpHrcno4VQIsHgpRY4nBFwhJQYjghUwQ0DCMdpspwel2ixa56p/b
0+Ph9A2uLU8mmeMGCO6lWoVdWBWOJf3hojiHPwBmjft1OrMy1QIRIAXW9jXDj9aGwNlsaz+a9kbj
elxgUMtj2Sn9UzWO592kq/5GocwPyhfnLXSAjFrBH4pgq8glkVrmBhQg5lkdBIvat7VYQzLAoFJq
9Ev3gz9YYRZmXOgjRIXxXlc0XrD+yLH9tVCy2HznSjESxoMGVniQEa14HklhcJI4fVzXa3ebzFKi
A9mVwW5MCn/Wwa0ykUwlXnO++LNA/Q1YAeagT8cezVk6aqbjTxYOBt2B9zQGzCZz2UnKZed4uaGX
7PhHjh7fMoxcbfthwuq9cQmlNMNG7FdyVs87NhLw+EEfxyM6mV2r5vYhoSxsQPt2gCmee7yk4ig9
7FOziBS7JfZJFGj0MUPMhuEedL3Cl8f4WZeT07ha2U+wDkwmM4Rx6jkj4Qh38PzjtLv5i3+N5M/I
VulZ7ZxP/j/yo0IdldjJX+b48Z78GXtIUsV7x/KuPjoJV8dIo1xjG7JNyNSF9vAMEvgqTq0hF32G
aIP9qi1abdLPpbNhxo2PDizU3K7awHIuPGE0UX09dnYS5ZL5Yh/Zf0jai4pUYqnGRV8Ns10ZlAaj
hW6Y133I5g9yXdEv0vJrXvu51H+IiXHQT8NwWQLb9YGFoQiEuujQ0x5w4wtdzIrwYLXn1u4AKU0z
bnGpREGm+bOvqXTKaMvJyBNnHpImLrRxQWrZSxDcZucGZ+l4wi5ZgeEYLgl7/A7+ynDKKH8yPj4q
I/nKdArgH9jqisiB1EsG44jethKpVuyrIBR+U/O2vg2nwEb2cqFhV9P4Jh0Jg3cCRP/2/Yc2aOQV
uRVd6x1YKquYmCM6HNlguvW7Kq35tpcM5pRA2zKSHIZknmhWYKe7oN4JJLCbHsSY7AOQ22/c1aBr
S1CFkU40UA+p80RZCPZ1OlxnwJEKOgmp6yn3/sd3xhHy5M4XKBr7uL8kXvbzUKOZEFMxDHyQD3SH
d5a4+0m3HVDP064NDsNoX2qDgnXT2wLfDPcGQBIfk8l3+Kb4AaB3ttTEjtp6CtYO6mTF3gxt3CEi
43nZUxdF02gkwv8U8DjZO/pfQywzdHvap0ucgKYbOssLkauiX/P6wQ4QvS2HFlWBuc2oOZOBU8i9
oRcgFU3+G5z8a7psLTFyTmSYCeEfHEGKkHkv3TkvEKhGs0slgfkXLkjz3BshqKq8Q+NhefUrRlBF
XLp94W+DxgKss+OxE/Ef0Ex44Jn/eLK05MCmuaZsQ3l1ruDtCmQOvXDA8w7wOr2uQO8QoI4xRaab
/bmCnORwgV8vIRxtg4cZ64Y/0mU2pyaSqIJk7quB/dqwPC4+32nCqjJaH0qkfCktKD4zdfU/ENav
V34tTSQNBj0YWZ+qXLZRb2RyQH1nnmWgvtaVIB4exiukKNAsllQ4bcLTkyxIL7EKNCDPUb5WAy7W
ZltZaWmJBtdev62Qy2k2GFhsJ8LWARHk+R1nMugaOSqBFvI3ElpCuKcOdPjVYeWC3mllbAad9de7
zGFDaOk/Mz9443pTNJGBY0ph+qXiez4QleT3FGj0a8WXjENTqSGCGIWk3fs9XOoaXWSkpF+kLLBL
M/pEdwcgbaJp6EzNly4sEHAhwnVwDkOEsYWqpWN7OEaD3P8gVEqNOh7dPZLmFTvdJk5zV7ZRopU6
uOZWxwW+cm8vWr0engX5wAP1lg07awJ9B9Yfzw1ksXnraiHYPuPZtnSoLSFoSzWBfk/3/rVEnBIb
9g5upYOys0TLmXqbMEW3ePjm643hiR1kwjpd4PLj/vpFwv3aIV0/y41tb6VCWyXxcYat1Yc2Gh4I
kFaHg/44OI4rIhL/yV3h1+2La/AUpMk8BZT+jlxmw61DEcyrqXSzusZATv8CvIh+9LH6DFwW3cdM
UtJf97DBBEyu1F0UYfn5+bdBePt1mOQ53Of9ofOuBc9LlWVDwwO6y7Pa3cLjBQeZCZ6DDpy1fI8R
5sxUtR3VyByNoPOdzWaGXNeoDOqWfSB/GDq1JVVok3NL5MPA7hScaqwPzhHaeFSlsGPVe05fP5xO
fjHXvNgAnRDZ2Tr3qPMjzzVHRWlkV+4Ihhjsyi+yuW75sYsq19ZKVJydIcLJ5pZ2LZdO6scUF3U1
wfAWkPS8P28AzL33WfkQNIFi3W414WtMBGYwRV7+/V8rO0TSqx/5C8B3c9ng2Zl/Njb16qNBfug4
OzYNH33PS/c5diHMplISkwa1mAtVkn8gzzrXNsJ5k4xzG5n5jtm2L+HKS8/1tU3VWBRgANV5+ViZ
kR87Wxp/tsWxhvAYptlVeeZQpt2W5oj1+UwRjQhaAWRv3l8BG5X4d7pRr9KcmJks1/0YLWK/ll0O
n96HC5ST/A0kGXxXmtPf9G9xpK9xMfnbJoew+XHIe9nMRSXIEbw6mrBvSvwPBB4Xl7vs5qLgcyPd
t06gsbDEhplaHTKyjIqAYaJO89wOg+RZlW3PDTgz8NaIhLrXGFu6wP8mn6o2HE6IwxBYzTF1nUSZ
xVx6fWk62mymh5Fd7NbBV9q4zk5ZRzQap1dfcLikpuLCO5cDwFz+MBeh6ndrJv9tPt40BGDtGjQI
o3dI5AaIOAa2pVK3LfPNE1p+FHxRTIt7LuO/wbOua/Bd430DjbnVBf4fkbg/Fj5E5JB4y4fdjp54
Jdeyb1CIN3BMMOfKMOx7SmA+5nkWgSOqxFkzr7h8cWlTrWLjeSqJwcLUwd8Uw1qwGglQ1eiwcg5i
uPdvOu+fBvQi1W70EP0/mQC7m0knZI1LlpCdQRD/sGWdaLWVxeMKIjbjgkvK4qAvrFlb7K7T2R1E
ttpZcRJLv9cnGkxv7XjBM/yIMURSXg7TvFN/eJwyGwqt6UDLf1mk6pqN1tCMfbYubPsBzHa7y3+E
ePS//BXfbO9LrqQNMBm+29/13XBOKz18Zn0szDQ1pNCVYRoSVDVo4kj92Z32JbvNhPtzcG67xxmo
KINqKCHj1r70VUQF29enoTzUtt/rXPpjuUy5QUl5o7lN9usCXK5whJ/qO0HJDhmWiqnjZTvLb5sW
rwKvs6Vgs5Pt21fmuMuJE6J3TP0d45xBvhvQOBOynSthm8GWd29nlLH/soNp64PJivmnVy8T7210
Lco86+c8J74U9iHO1rQ9WBF4ucMmUf/4GH9qo3DktoLiSU0BtSvRxJJ3s+RGnbTDkRFaV7OE5awX
5M5s1DwJWk0BH6v+JPdirubGQV3HshF0h9flIpO9wgPEvhPyVJYE+7s6zn6iSYlA2rmIWY13/Wiz
OjlOgWVk4SDL5gGiLh4ArwBu5frqVgP9abNpg1GmGW0aiJk5eZ2TABckR8wgN402NCvRNQ96nyIv
F1xeMMDbft61He4o66twZWk0tcwh/hOTzQjzKUf1hppQ12WBLRLDbZEi4O+64n5AJ2OROEnFQcqv
GJ8i54a8yHNOKIAsBzkhG+azM6WSL/A2PHbTQnxlljlDanWWytCHQpmprAys/tf6tv1tWVs+OUTc
cOCA46Yg4PnCDEkdo667aEAbJfYuk1mBx1AY2sQDSIIBnd++ZSrdU/uLCxtjMtPbPNqlJlI7Nhot
ihZjy6C1hezXpaduWUTWUvao5F3wHsXcwb8xj50GyN2QcAD2HfLqp8WNyjDv8Nl2AQcdQrydz6n4
7rReKuDp0Z+jXpJvsygP9slnChqKDZazQHtfh1oafNtMRbBbf7RGZ2Sl4ZCpLn5olfOZ+hZwVQxo
wmGwXmggKbifJS/GVz0vsUsyqq6d7L6B5TuuysihViq1PGWpOnhpJiaGnmuERuOaFgjGth2sXNx0
VJ6DwBJHb4oU/fFGc0glEd/C/wiiK4UYIHZgjocrIxo+xH9BySkE6nOKufXVp/LMMrFU8F8oFfPv
80dXnsCuTZttxKF0WJ3ELRATgkNTQtAK5F2UjZN98kTyEmMD444cAX6hMK5h/wUdFQCEQJbx3Bn8
jCaKj7bjdR+YM5PcIWHOAEXQwRPMGYnL96TCD+KcG5E5NtllXx72jkgOALM08PkTi/GQoFPnqJFO
rC56Wz1H8B8ooSmeEv9hq0crVsQGZRi/NiG684xQXVlqQ/cAlZovvckh/yZVwnEk1JBC2t/TvjEt
dzmDPN/8Fea96Tn6HEXcd/6CIggkfn/NbypJ6H+JVcD8pINx8gsiwIVJLXvg49IGKMyk3pt382fB
26KPtupIW5RFkfclZZCK2q0Dhk+QS8USsJSocjXLoHp8YY62YIzMYfIY834bISwTfj6S6xhxgSUN
KSZsuHm0490rAOr5vUzwO/hae2UZZJho5jckRJnQMiV3qBuiri7bMeM0TfFL+n+kcY+9OzartH0u
lqIvuLkxE5ea6cMFwG4pE0r0wsyNnTgNygU+wDdI4XKuSB6PclgElCPJjX3LsF81Gm24EMBWQpb5
1VdqSsQvQj/fwYIdobg60I0PgUBtAZYO9xNxW5Mqt4C/eg1VR35HkK+q0fir5yEipMI0m/JzRvPI
8o0XV4OVsi2O+iQoOlw51bKlI32JTDGbDapDNqD3K4meRc0jfYPPDdAnnIbZbT6MAmwIpnxwHu5G
DnHohcIicEu4Fs293+lP9pBD4DUWh6U+J6N4J+iqytzRhM+R4MLcuFbFmdfVhdgwy2kFDsQ2Q19g
8FIdisOLlQjO+mciJc0d21CVy0SnIRM3If/GovALzwBSzKBwURiDAJR/jS7Oo8YgdlTOOgxw/a/y
s+BcfNCP2luR7sIUPWlk9QOjmT+pL/C50iigNPuOTbq6sMyy1poFehlOdmEAJLDyoWXuH9+CI9zC
cHV5LvhCk0VrNfTyCUA9KvsLSZ5R323yA+nnt0G5NvEFEuxL3Pt/4V9qgrIQj0Ap4cyxxP4duV32
kkHlFkcQTRb/DfcL4mgKbfShN66ihwvWZD0Rn5AWvRtR6XuR/6Ql74gT7S5VfWvf6sMJzZVPuVQE
G/8izpED04UtgbK9TduiDEyxF9V/Vs3R045FOH36FFXEnrMe3UrVGBxpQ+jlBB0IoJB3nP6zJw2M
OmsBY3ZfxENAG9Drnh3+cWYr96gNnz5P4NSSe6gb0B5h24yfzivC1C/h5vB3PJ8xp+IhPhtCZOkH
UWL31GFve9GrhCPnBtygR9RalSwk1XZXdQAr80tsPAiwV2hOs1EkfAUmNM05/Z/QSuEdXRbO9jpJ
LkzosAi7IpxvUn3r/bOY7Xq2ppNdIorswNepyWB7G/DR3T35hM75qbXshD/f8TCdgZjME7mYRbyv
sx3NvgiNNFCJRz3FuGINqQUxe3KghYlknnee0FUjKk0M93eVDoxK5gmMoNQJc133gcC/lczN/YpJ
TrNFXLU8IHUaeYoQbftYHdc68w/hx/5+uqbhz0k1/aPZXf7NQTMduwstD3Q36sEi27ijk7BY+bWP
qf9G+7gxDi2jrYGASxoGPWCyBxz80wSa9lXyx4yaEfZF/G6eTY6gDK6G/9sjAVNc6Eyj6BR7WGN5
SBWmsKKvkR0b6rfHyEQRQqxxUjM51yxjHs+PwY8Q5UUevitz8meESwObNwry18/4bL40UdAAbn7a
ixqChE20fooymXw4ZlWkJzjfCh2edC+J/7o6N5TX1I/2ArUuLuDbjlBiaqgi+gjA/XB8WI2zKCFA
FQPrvmsnWEQTA8pxdQFfa9hq6QLuYR/APjhgVjuuaWUcDDipoIEs9OBvgdIDsvxX3kyDFlr4vdiv
kvUm4iuKKVq1EP+13OIEB8zMxeIANAGFjbzAWDPia2ECSnt29XhK+M7UU5sWKLYt/dUTeL9usfhB
buhfC159txYR+cUR9CLCT68gbgm2meadezmlTm5rcH0ShLdZjKdZ7td7KGyW1t8Ek1kAER4r8hVi
NUrj/UnWdwB3BiW/HCTsiuueXUD7sKCOTjpRhPlfFxO7/cZCORFhhUKdvU3gTdS+PVyW45v+ACMK
TOo+RY8qURPna5VtdnHgUBjJqo0mQXJ/ccWWSsBQX2804hhBDyyVFPqbfpCLTOOhpRY2LATYiSo/
zA+QXLjDbSoAh7pOf8WB5dgrVE7xO3qkHG1fDDyOFOQm5RNJNw9idF/3udluq89qde10N5yyAz3u
rCvhuO6xO9XFYN8niBySJpuRLD9JL+CLSYxsNiKzRAcs0/goRw+AUDuvqicI2BhOkXrhluV2xi6s
RqdZMUXkQqFqt/90Jf4YXrYArTKuEdNOKwOVPxwagZvRkOgxn6o/yiHqAacDUS9fUgJpOSRqeZ4q
skDYh3FGVQDjyKqB+y+qVsUoJ+w6A7B/+ezJsmOAARngGLhURbp5RMx3xF03GFQ8LC2iZ09AlPfX
Ct3UCAzZ8jwBtrKM1YFUgpitRiNpj+yQpjXdB+pJwqWXPaV9rpB26k6xHOXzCp/SrhRIIM2aImam
jh1A5bu7uhw3n11KTNAihS6Oof3waiW5kbnMLWnNFt1QHJJHzGslipPCPhyvH1pE4BuBG/E8tDyB
OnziHC7GLy69hNdFMKIt89zAHH1TwM0KfoKw1VU3XXSpt7yNFQSjllCF5UtEDd2OLY9LeiYcRrK6
rnTbzJd/E/hRMNH+c7TCZG/BTbBPKp9vj5lVtMs+m1fyGibC0OXv4eupeLrTVdFaWHw2nqmWjEVn
moqSeMZfptkDOYdPmlcCt4esZuONRS/t2SvX19+PYZv7GR2tgwZLiplr8Sx1ASb9ce+C/GfUVRRi
G2v1z1vUVD9LtmNeXgLIwred74PB8l5lzaRI6E+7kP5JkxU/mj0rxhRd6+lAPBFdux7WmuMzH1Qw
27/H9ZE7jNH6nODkMT1prR6usY6O9102TlLWjpFNK/rgtsxp3l4/M9pjPW0ftOY4ZaRxXr/ByzLh
2EK7yT6dInzdeOnWR7emGAxgzHdOoczTjHoaiYY7J6TnY3ASxgUOPQAGg4Xwc/dC9lxWIiEg0sLG
yWji59v4Ep/Jr8zNeHU35y80WzlqJyAJrlNqF/0oLOyTSaj64Wfl+0XIWNQOPjMt+fq8r2KIbkRb
doFg2olb3g/vub0YXH6AcoBRpDfhNnYVKdgdHnCqfwN+fIUrji5zlVyuDCZQhuZmh8RZu0A7BPtV
kdE6DgGY6hEQNGIfkIfb42HSDZs95wPGfS7vGGIJ++M2o9mOxahN1806Kq8mDObLYi969Ubsi9tn
a2JED9EXFnn0eFa/FNjUjdLeDxFM/qOjgwpcpCckaztW0K8VM3Pi4Y+JPo5VNKiFAJ1YrovqT4Ww
lQSR+UJmMxQPC+ZI4hLqqLgL5eFB87tmE7xwxQb5e5M9GJVzOoHIDI7i9XNY7OvS3CXNhTgL9Ng2
Dug+d+EiNf8FUVuLdD8dMfH3mpZSfwcThVETt2oFHucK4Jt3FaHe7FVeZ+vPgBDgQ4nX3R7GKgNi
05KBJk0iVCnSjdNZh0ZRtzrhmu9p1xDKVlOL53qsji4TRjoXKggyb9DcNGhGJ3aHieJ/XzT/1d8Z
OJceBMd9mb4h2nq+3hmiIQudUNRuaXNTEWczvyJroqu/334mZG0wO/7IyV6OSuHbzB0Rc8Bgy4nz
P5DyUmhWUdAU4hd4R7gdszafGzK8X/iy2NGiED/w5ATPJO2DTnY2XXMkyxXXh4RY+W03rZFhmxdR
3XLSLFB3AXwpcavkW4U6M0fruE7rQvTkP3NcXoXFduG0jc2dixV+cTX5rHda927ANGd0KL6Y2kFG
xjDw0no3FL1aRSQBwSAefDTNFKwFe+MhAtqwFvdbiZh9IikXSmCUZxZNd99ipzN6rgZYJePibWIR
T1sOm20GI84cYrctAxkIQhQssKRMYWwMrHfP/jVQ4UUKtICGb7YpZ6gO+ujAdmliq2AhRtyxanEm
4KsnfhTyG3TWLx3EHkkJzZM4P0mOPHuXqbqmUMIGpaBa37u9XWV0LJU89tJR2a9KeKdMeYgRxfdt
uGH3FmZPZ/lOYHcRev9u37nP5lkz3WqZaMN59CNoxHUwfHtEa/nqep7SGZHKVZQODqRFtdNL7Ijt
mItWuJ8zPbqy8c8HKfjtULehzGoqqGN05ukwFbkYbMLwg0DicUbicGZHu/o5JnSv0qII4FrfhQr0
lVaMqCbOcbAfT77m9lq7q0ywm4VuHYAHSOvTGfOQ0zWCMnHnMIMIYEsxRlRplvB6obfO7pcQiYl2
/r3yxuuZjEWVv/3c8AzHhjomHHz6lxGeWjp4++iJDUi+RJ2j3ePaAQya78mn1gMJ8t4f3SG4H4oV
lD91t3lZ2PM+QVJfFxQpuX6buXTAe75g01/kXOHSHEKf+JmTqjB0DZdroUN/dryAx7Nu8CPwbldD
FdsSTTKsemYtPC0U/BP0gfy4w4H2kk6oE3UF4c2xyawiRxUMRnbXOvO2wng88MRfq2OOpRMeyFZD
NHgwYC6fkix5N0VR+0lxLzohyM0XzaNRDKJIsjIcAW9rdkKaN8WBAt4RHoUbt2nGLy8TLe7BLqAE
KAZRSESbew+Y2DjB+avmXDaQpwV8VibFT1y3t2C2rgpAWmiEx7vqu91NyZ2iax+e2EX/H9eJrwSd
INbPEQ/OJQZbozbiOfLYgpa6aMlom4iin8MCaX1bklF9vc9zbOwDJ5ehBviBgCbwvc2Hc3RESlXB
3PFHw1OqPG2w83fsXjhp7J59t+caSpAu5wdYE3qyCRTvNbyoQR2j2ggKTBL3iD4VG/1FXIf8N/vl
JCjFuIfGL2FhQQpC3qNxXqj2PD1STmJnAnbXgpmzfbC9ZL9WHaTJ3G4UJpguc/3CC4gvHobaAJ2e
OluSD6WH2vOMCf0502w9e9Zcnci8b+8b6T8V8HeTsWTRty2lNA524phVHx/EN55blaxL8fC/+1H/
Tsy5qPSW+4esx1lMCaxH5fW1qoiNP2ND1RAL07KURyXSGYTKeGW+bVzJPnmls8rx7C4wYMEbqgce
eE9FafDehjczEoIkK/o1dW+CajNl/IvrMU0tXsDV87qGbyYu/lk8KPa9bxVQS7CR4Y+QS3DEWdhG
M0jZbHaXtA8Vgn3/UYsCYJnl9O+E0yzVO7KXCRxRM96xBWEK02Q3kp9MqAUpjDbG4IEOHr21XE15
2c7B7BdlJXVXRDbowNmiErfF1FCaTvyPJ4v9b8jMI3Nz5Gf6yeap/B5cbnP0W1HyD4FrJEzFHHwm
OUoEYwynURoeUi0OGBDxnSTSB3VTQNgOkrDUiLf31LcmrKzVXtbHGd3wSnkHqhXe/FVMhnjN9h6l
O1Cl6SQFjRUiYYrHIYRvLI9XSbTHn43kzAoKkDpvIDqHeZmGGdTfYr47dRDgDVHG5IVYAneXlEYA
VgzI6kEUJ1RTvRk8Bx4uIJ/2YT1WWOCq0h7nzzVKM/oGBaLjMXh/7iVb9/bfjL2OgavhDYFv5du2
3eo4LVoJmLH9T8dZ1W58H9pgL8cEfupH+6y+SGL9W1yUdLJ0yHMKyqlfPCwushnhIngcIJvrN3eO
tljMrBSw73823VaHhj8kD6XLq5a4y6WN++0rNnWiwEOHfrP3NWgdBfe0V9Nt09j81nxCaXlLwV8g
TnABrqi9W1bArBXKVe0CCFBPKJJHgk0opv9rwffPtf4syylMSTXNF6Q3LDATHlUnb5Uvr7k5yZxl
O3X0LqbJLmNjklSgUSLRC/csdCrF5L21HVyEtbGzKcSDqCLMSHTwnEtMOshAYuUQjUT9yQD990mu
NiCksKPDfaVLV/p3xoxMRzVKzzMsSU9uHbR4f5QKbSvLe2RYfGY1hli2nxA0OsatEaEoDx4PPjfj
DvG2BaJjIV/JnyC2vSIZ+fY1H4RvMYplzmhYqHxooJ0AZH4E5MNdoWk422mk4kr6C9vqOFOwoYSZ
LPQec3cHUAmQ4S7FA6dCuzll07vzx+6lTsB0kaUmN5RH9+Xg4lUwZ4Xqc2gRQYIdZrufJXtKKlLB
QA33YmaYOCSSJFnRSHR86jZ7DHSUQjYajyUX7fwjcu4ye+Mbz2IYeRF1P/RgddPwaf0Lodjh3sQE
QRxOkEYI46gbnnZPzM85whK/4g0YpjOmq0zVEsxdGIcqJfWCRFjopQvUXn44wlrhWI5l8g7sRTFY
wlGno09bODKYtegplU8OO6WdtkwcImYagYfC3lKrO3L0eZeMJsmvn+hj8TVtkwMU0EtRBA7yZPIa
/u1gxhjvMw2riGOV8b9GoLmlaJ9MSZwqRs91pa5Qk2pGezmzyKu6wd/W2aRPmcCx192hxwJkBhvw
5b9RFX4IwcXK5AZboVITUEQmaKGyp4l0SjwBFmOpkXVm1wUqCV7WFeXvh6PwvmxC9KCylVAhc1f0
vs0EUysM+EeTFJjmC10WlFyCsKvI2zySPNVFa+hJlPvB1zjVIGjTPiod5YJ5wr1UDHBuplLJTAGR
O5wMbdxW0+j3V/KrL9iYl3Ar4y6LSpL9xzn5b/mRH89VQDcrsMEsGBppdDpoHrNGoRdbJS6IF4yH
DSCpCG8qCnDCgFeftpAvkCHI5aBRrhfjYRMMPh+dJA1zEth4G8iZTCCHdD2SzsGzw5CPQXXiS+EV
vUhVSkrZoNdmrEqXH9buvEVjB3o4zy5mHhNvVoEGdZEBOCvdC7dssD2NG9+azlys5lqs2NXzkFrH
AEEOii6/xcD09TZqvar7yZ4R0WQlQg2isVj/y1GcOk8OXqosBfwCW8y2R+ANxWBdwrw1s/NqpFul
PNlAULBrnoxYsaQG/jO8Pcps2rxbGaxhkZgQ7DofdU9MM0KjIxMdlw/dF2pNdJdb1dYBqXi4x11I
8eIao5a9Df55VU3mBKG+J2jPfa69AP/H8jP+Q6lKkpMbAn2kG/bEkKqDdg0TvmYv1M9G7vCAXZIw
QwaYfZoA2kibwiV+xoqveoo0ukFGSRHMqyM5fcVADt722QgZ1efb6O/ai1olueShNioa+ZUnXFCX
tQ6e3r5Y3vJcJPprL+K6l8JS7hAJb/JXkRASVcx/aWfNsPK3AWdTZ6rV/G+u6AJUpGvV6gd8CYt/
U++13L4ST1TCEAQy7Ryligo982J1DRC5CPmXfsSUNFcnxYCaL0GunIFjn83niV7As+VC95mvamx+
158Y90bkp8XiTT6aXsaV10vaQ6yNsht9+vwX9ALcALW21PplDG42Tx58ewl5nPD2O62geDiHE3cf
TxufA8bzeCS1HSGHOfZXK+gWf2+q2jSjzDyMZOi3U30EeqVx2TrXOvRKDLdghLz7s+ZmEqiKV5to
QpPpaLXnXmeu69w2qexNBqEvrFkXfnWAmVw9dGW6Auk2gzNp9Eda1YbPwvijzgzv6akgMgBE8l+r
dqdiC0pt0FuPE8sh5MVKvpU3TIdVOVt5MjOsbJ9b1hdu9irCPFShbjQdLm4MIPlrwGLGKHkuWocY
JKMSngz91AIhN2wIzEyzYyjTy9prLo/WAokLpa0G9u3D3dIo7RCPF0yMMjvsxARkOcmG6DA7orAF
x8wQ6qa+TZMBaDLEA4/eBQYONndSvSg2QIfrQVnXqp0v73vNIdQpnTgVsmv8FjfWM/zYH08QczUw
FkXeBK5b8Z0I7D929a3NJv6BcOpPxPJIPCOgRqrpJBKGUYE966x7/H4bJrrCup9LY1X044IvDBrw
QB1zLJlMHeYGYk4+VcotvzyX70hKViNn91ow6c80oRBi5o2VR2BTS2DfiDh3tdW7PzX5+SjyLkZj
m3Hvkc3KVff9li8NwJKm9pO2AgNZDQJHh/9LAZ6ME8okFmscFqH9jvTP3zLg6AXvz1wnyYPcKMIO
M8awZ2kjnYhUPpM3ruPeFtTYlw/T5haCZQFppB+AscwAQdJ1ETe22+xzbKLR+I2mki3fZHtqKVYq
aWjBD5Lspve6qI0TGN2nx826p2VbHtAIvM58+crE5DQsFXT3v1wzocf7NL0PmN47xspUWpRwBP6o
0u40hCvh4+tf6iOpVAecO/XsCrytBLPqWzn2Kx0ygAecL0ZzZxhKeTiwbqXb2ElSpTTlu19z16B1
PzsWwsfB1vsx2qxIhgYVDFSV4KQ536v2RUPKDx2leaw55WufJFek2NzFCBlIvoEQLeRcKrcgVb+x
lUH12aephE+lHRisOWXgi1ruKLp8sutD7lb8Ufo5otiXFw1sNvcStLVWG0f6kHlYxTDqF7RVg9Pn
9TTn6g8v1e2X9DYCbGUyQRcPuZfRxFbqQW59cj5fGjO6kY+zTzOXEnhRDIGOEDA/I0NCM6GUpbC6
uVsdeVMkGvPTGAYz+/iYJCWkEBc0jULniDLieMOYMx1bqsmX7IjXWpPRj/vzSGqG5dtz8RRQkrzw
CafMObJmC4kam9KogxvvZ4PMg8MeNNrqvoBQKLSCCOQMwCX+ROuoxluGOaY+D1ONLN6S2NBKtXCW
5jaLsFzoCak4KhY20OB98nOq9e9up4xuHH+J2vi/7Z3ITF+hp3Cm/m43123wKdl3EVVbLYbl+rOr
dFLx1cev//uX/cqcoXO+2B7MjX53IpJTLh+RGkGrFBXKVQvYeiDDfuD/u3RKAIBR/YrsDUjn8eky
2RTfkqSPIi7A0AfH9IHKFqq20d3OuOHmUaU1+Zn9C48nlm6g13AaoGGBn6jT2txgT/NMuiiE0nY2
fMO9WYwHHpagIo63vuTb0YJicd6DPgkTc5nT6rX8Kmg6Hz8Je37YbnxEfCS/qwPfIyER9Z8TGrXZ
kdN0sgkxQmRHkMP2SGDRh9xxTgZP7cVYDZPk44xD65ONy8ZIwauS3JQez/s2za+6cTmnTmQGcSz0
i5YTr8fI+QwqV2USHYWK/TD8mGMYdV7WtZnplUH31xCo7u/+XDeoKFrN99CBgNdHDWNz6AfciC2F
PUMnqKfXUxTX6DKT1zbjJodc0T9r0CzrJGQwT3pVlT5eNHhpjdhkkq8QuF/ft+EXGcMJEBmT7zX6
FBKPL7Rk6ndMW/bI63lXyt0sXCiCmWOOCA8t2+R9uCGJ7xT28wzlfTRNHV3P5Jq3iadtYNWAeOit
Y4ntTQvqBvaiXWyBPPaYIWlsuNGrilULLqODMKiozlO5NQfHFZpCDoVD34M01gaac9CpDNPf+jM8
DQ5DGdwo08fhcbybxuiKzp+PrJuTordyUHyUqAqBkm7/JJh3lt4KPxHODv51ztQgA4ahvywzs1bq
sR4y0tAqyCi+4n+79yQd9b5lXDjB4JH/hIimUgwVd3k+Fbumf7QRBnOlx4Lcat7OB28an8aqQQ+n
m6i9yoMfo7YpFqCBtw1g6xLO5161jGN1GrfnkTOCnIqwSKzU+nkT43+AePGQO8VAobyu7nQgCbIh
PrLp8B4JJQDft9wc9yg5ZtSMlkgbaRzdrsRi+SMDabwwZY9UPKojiYgERZtrZ8/UaGeYtiGjAp1v
82C6RwppJdScx13QePr1ZEx47Xz1P2brH60m6w/OIvQmHUN0py+n6h9tSD04N5lhqzGD/+2NXPPG
kCyEJ7LqGezz3uJqpgIJ5bxcyGVj4LIEcqK0nTRyFhlg+V8BAxgstNT9/WHnxx7i6MdE0apZftl/
PiYZrupAwluyLUIjfV2BAPAIZvBeLaGLHczysGUnMFjFrfq7BZeMwLnM/LVNzLE7ZWFhfx6Gg+zI
kA6UCOBhLmsohyAmXMh1coFRob9KZnDGqjUCyokVpwhczg2f1CcjmXXcSdWL8oFs2Bkg+xuyRWBy
AiHbJulXFfIERT7TUsTh82jEcJVaXvEmogwZ+du3br4X64059teYBmchtuTKivCc5BirKe+i79dD
zRlpMEl2M/zmuOxgl4igYo7cPYI1j/NcfXA/HTzAmDH6oLhMxTaFq4mhKk8GA+4XkaDk/I4tkzEX
eCLVdsU+NRYm5aaRvytpw7jZFHDAlPX9AFC1B9AW4uU/mFEBt3vThQjQLxzMZ3MzNL9wA6doaT1f
59VqlFeCNfhQ2vIcGCDb2jO0XN93aQIjWDSjQ66gfS9zkXkzcMt6dvx6w2U0VnUFkCgwZxmf/ZU8
TcnkFEIE33luwMA1zlAi7H2aGE2Ub8XM8/hqsKghZYTvPyyOIKuOChN+xxpY5YkI3IiYDzbeFVN4
NWYOk/Cqp0tArW6qserNEyS73N3bdF4uigCkIswf4jUR1gqhRTmdp1KUfu8qSs77XV4B0773Sojb
0bnllr+LRVZ0sEC8yKEzFv9qviQDGfkw9dup5Y0KqSFGHs0Aqw3ag6wlkOJD8JVF0dfsoQK9M0F8
3i+dLd8is1dj12Q5mCnWv0I8dCeZuOraZu0Tz5dSF+dAm0fLZIgyfsLBRAPhSnLR8y91ev1Ac++u
g8VgdL/vFDGY4xbhTmzGkIN+uZvbP3BTIMIYPsU3d/KH2V/VhIaRaFsONVCFz7yqdsw6NqqmcUQf
qRCSEQwlGwSVaJJdBZQQ6atFjFcXr2O0DX7n/WG/wSWgYalSdJc/jrxGE0ODJFH4mgSVFMhPeOrj
N3yk24bUkS09Vw2SJwbujpzKPbH8OW1dhrMRDFJCbuEM+u/gkbM82LWFym2yd9esAhy3ywG2B7SD
h087XCk7q08iqbZoesTJLa3FVhb5KotTngNqBmpMFa50yGHF9FBlHcuXpx1y6hLqWxhQYb4cNz3O
KMsT5Q4YSwweW89LXrZHAb8HKzzkoYIA9mqFPkvWQ+BnfVpV3ZxJ/Hl0yzz1RnB/qeArhHTp00m4
vbs8Ch9zOmbh085O8WfvIRlmqbjFwUgDpYd2zsYAmjWUs3RtPCV0V+wOqdzqvPLH3pOPXruaRZQI
Cy54vmuLV+0+CMesXv1M4at25kC6uNZg3DiKZCnFb/gi07h9SnQI8oqKgR78rFOUtIymMRFfBUu/
FiDGxyyFhdbyGFvcJjuX7vk2ySj52BZIkwqmi00FO4yuN1wnQNslktZPkK6Fzzw8Sg2RCOLcEd91
b7DLvI9/uTmWRrzDx2KhNrChO4EoxFpw+uNXvZw0BsiaFd27rkiuy5u8aYeIvQSacXPOmmjJR9Us
YizNy01oCOulb7w0WpIcJ72FzgD00HBSfJGOLKYRzL9Eml74WNv0mU9INMGpoRwXIXh5DZcbdwXq
ydcphdjE5BUAC3OdTYyRvuhtrdIf0FAM0HXMDMfONCUcEX3FYTmpVFMvuELl9kWrMJi/atCQ2aaC
9VyBOCmEYyohkbYWMafu5+YP+8KFCLJrjWc2XvNN8aXC8nzy4REnCslRCbNqb6sgz3yn6JUh4t+R
EKW8vrthUvvv0+Aake8tgXFMgq4qTXXVXBXeea2WjSGyFnEVyXw0IxOaEdS01soR0dsb8UyQltFD
gK1j1hPajP7sLCHh9uUf9UtbZ6q32kjKIio48D/mIKs76Ndjj5QHREnBrEkQNQYdrvSo/A+bzyiL
e53MROc7zmMbWT3eBb8ya9qDkLJ60WFyttMhgvvopRt6f+aM52IfsYdYv6GSiBkr9/ShhIsWEdEA
fT0TTrThV6Awifs0RuKAMa9l0m00oMGMnawOKCviVXsGKAnOpXRwuCtN0YywQ36Dz4qQ0oDKr+f0
y+pkp57ngyW525x8KSb9YeSBu33WZdXBq2sOjZzaKabR8rACVa0TcSoXl80HXhqqmFMV6tvU21IH
sYLctkiG+FrqgGUOmbx34Yg5MNHXEFrF+VWS6N30P9VAa/uisDGY4Tkr2UOa+r8dvZ7KTP3lWDQ4
qawI8jxMttmLftKY6AiYyGU+vmU8Vw/8FA7AN1PkvKUYV6n1mG4yEe6oSghOCYFgvGZ+hVCCnzLq
rhbVMLgPjA7h5M7oc7Qf23/CM/+CjmOMQ8BBN4B/XfuHtlhdBUNTdIzJoc5ClN7ue28l3d7cUFm/
9wJl/cqO76LC0Z4kA4f+scTmNOouBed7ZZpRQRR9ct7ilWTfDL1xj182+PpXSlBnacbULOWUW4cE
Dj88ovap2REL8rnMtpINzCR3LC3s/Leu1aE229Pt0OWk9EwriVa00gjlB7azsTYx6VMdMwkX7tY7
M4mkKBWx3hDqGOhs/GAQMmv7sAqAQb119UoyFs+RqjLSLrYiHeYOfOl+5sD+jKplP0AKrpaZ4xMy
IOBRLREqM9pJI0zckC2egeRUGZC0D/f6ffpLcSii+A27rVl8HA4pEyMuaj1xqYsO/PbcQyxLPH5j
sUDEgZKaXXRJ/+yWYAXXXAubtZulOfspC8B84eEqeV4uuMliL/aHrS7nCENC6LgEUA8bbowJcpzM
KQp/1uECXqiZoqJtUV7Ry70UBLSjKUneiUApKb/dtNJ2ZuFsYGndpQqTNCnFx3icb14WGD7Ev5LF
SmLn7q5cBO4f+zffJHUcSUvLJkurWNVwtU10D/7tGR5+bGiujyG08yPciIkzl35SSyCW0nmhVNt7
gmD+97ifuf1CiW1RwJk7OHTQYjKOKf0ZmbBLqr8gGAYTH/MbiGteovJYEFFHQ7NLbwT79RvUpKRm
ctUo+GkPgRK/D1Nm1QnEBb9Zz6BuuVxO2GC8dSyrpI/5OCzToFOFrSdwdShNRp+fLU/rRAANMrPk
43RNMStJXRISnaUyE4uHHb3OiEq+Io581vFK8/2pZ99qAolKBSiYQBefoU0N+SeR1wMlcLRyGrxe
F6+naFRctdNGQS1wflFv6f4Gx8jY/7X1UvWTM14vRWPWoDcGyB1WnPxbhAHCJ4DxCha3eGC7KWiq
7q7eM4vdFqbkz195/1v2TGt+L9BZF+SOMhQmxxB0mlOIGvt5Ug30QrZkXFV0lSb1WoF8VWsV5xic
jPeALPoKsaU7lxAVKO5PrpoeAuScI1a5sW36CsFetCmNbzKc61XcfvxHmx8Cvv+7eLWDdGdSQhkS
0u2dyEyXWm985eV9xac6fRgxDqt8LXpKd/oIFUuCnB4ljyDVwVwOR8wj/L/yU0aV+CloslDREJee
xp/Ci04yJSoog59Q4ejq+ybc2dWu06NVz2ZwxVAgA49QD++/HxAiY6PwBL8B2Flw7hzMeHBmpnCS
qLUvuDgK1mn3B2qZZUV/VE5HaLgqCzz6/1oZgUWmuMnMBMz4vHlGE4sSLr7Kx0Ycp6t0+gq1xU/Q
vRUALy7HE/YeRnU7+49XlymkECHnuYgh3KDhaLpJSTXRbinQZstyCRUaYkmbtvzCl3osQyC2UcHx
3x/Fx7URNOvFE88jenGTYWM0fXFN5ZDVhNrJccZWcUEbrwwMY9NdePmeJLnsW0d08ESguaLIGPpc
0qt5Rehxj62s5+0QWRoZtkLyuB4J/nTclDK5riCgaxBLVPNc6Zz6jj+iWxPmQzJYPKGOCe+HRWWv
vh63tqC4Plvqq8tGWREkPP8chVhj4PdTyQ0QtYFSFd5CVqUHzT8hJ9Ltt3EL9wih4YS9/l8ZYPRR
vVDgv8nftyMxQ+wDB0N0vZy2tZskoHkR+ybNNJ5Zt4wOdMm1NebI6AmINpzBQ0PYR3rWWasonGaR
udPZazA6O/6dIKokfBSgLbVzCCpVRvMNQmewYTmCsJfiNyv4kWzW1mmdB8qcnpYfVLzjyeXGUL0k
v90X9WidE0ZVmGQ0zXj+bY7tq/Xiuy2MRcZkOO+cJkI4KdQSBBOv/ahXhCJz2AO868plf4JHFzFB
Q8qi9yI7lmMQEh/Zyo2FwiyGVuJPAbnIv8/0G9IEVw3W+PWRA8MjzF+VOtiFQ+Xw6Ulq7dC+4TIm
bQer6/XKpF7XYVTuQgH8SrqSqFk2sqzoKz/2c3scNqVXuDWfHD46iG9Ndtk5Q5wMhh+dHSk+TYMa
6c4lvJSe+PK9SSqgkW+RkHZfYSZ+t+s1YscBzL+JS7/fwOBmzSJ2wC10AIPs8LPRIw6qrfl+Zjqv
NJ8Q1/S1Uvh4HHFysY9MZ7XT8s+v+gkRqYLSRcrAMHzZzftTFULnmQlTIFhRpveX47/j6QEVj6gn
nKsqJRg7JUjHPYziYPn/C6fN2rqGMAah44cy+C/2XZ8jJU2WjDV1YE4pQlNA5z1OTZHn38+NMQkl
ikdkuywW6TSQMD7OBoWo3E4rmn1O+AilmZxHIrpWQ466VZFP5Z1k9urDJzzVZ/3/h0VGCVlPvhK2
/073oMdYEMKlo1j5PLcLmfUxBgbT7BHLSgGHjPKc/tziX3DHk6+wtyF1QMhcV0IVh/BPoM0fQYSh
xkx1PfV1fB/dpSvrczIr/VZDNk6/dtqncQRBtReYngFY2nl96khFFCr6qYmRpN+8+yFm+pyEIMSn
B+03iOStf/Qk17/oSFCT8thEnHNz35QCp4Ej//eEjlFU9SDbR+GJtiPFJDxmEmzncf/QDtPwXfIc
DZtnu6OQKIPLqQU9jIAZ8c52f1e2V/ALi57mp5ZA9mgtbkcY7723CYNkpZ1Bgede0oxdyIRFTo09
6t58rDh0exutelCHneY6aIWa1E1Itoyz1zLY95CdwOGdq++ZmaTvcbPYU1P83vGuKWL5/lTJGphA
nhBM4UbfnzPtnI81gnPzi1olkdFlrQ0Vnq9s3MG7QVBQL8XbgyCRNqUnrad14qn2d9D4lJ2QfxK7
lkXpvyl5GNl4KClrNtdTFsNMmbnK1hAKKQy6kCD4UwLjh50cVAeyjrez7mBCwUrxVx5/HQwnfcLD
28IrCSEDo0Ej360V5YSUApIEYDyysD4iZAATXio96UdRN7PPtkSvCoeATFiVHT5lEBguUhjKwsZM
c5ba3q+0697pfl1I5oJBYlL67YiLkDJ6/+9Qha92LtYDIVc8aELTtDW+MvgVH/STODoP3TTmAC50
apBNxeZRMaxzRo4V4QAqR7cwQJ/ob+w91rkAIJNcS1HKV4Ps62tWYNHqPhSWLFn2lKeHdruJF2Z3
qb4zSmwOErlvHp6sisCyOS2uSCNzhvuoZMHIb0iQXp9zofPSJXa08wkONDSkLkQPwnGKZuo0b+JF
Qp8QhWtEetO5qQZDO5vlfZ3nRWYMIwUcvTj1KnHEVlilu0LVHjZU8bj4/7vlGZg2LmE+aLvHhtPg
TjzXaUM0GO55bngOEa7tZUxg3mGFlhQm+MU2WtfUhssPzGGeLm4cAkiIfImIa7ciTMzaUVxj8kJY
DmIIoBcMN91qmJMU+s5D0f8jqpYBLrjIZqhTX/VPukF5y0mbH0cxNb1+KYoLzP8SJwhq7/W4mZfQ
NvfQRY6yYBpbbrHJwobUhiCM++EL9lm87rpaEcm+dU6EZRaHm9KWP7rwez/bY6NTMiuLtqJd0UG6
NIMffg0BxSAJB+OZ9QmenB5Kq6//JPbr678tp9qmm1CKuweTfiuwlUP2Yc+hyqT6I1hTE+5xthQ1
tB8vl1ZgwfxQQJGvrZxfxlvh74Gye9u5rczGZWPqsFj8cu5uMY855Pvlj8UDRO7MD7aPeWvURPLY
FvFaYcBK4xm+0jKC/+utPa3342Z5aMOiaPAW8Cj4a/2FtT/hXbUCaSVMFIhlida6MK5fZMRW90zG
I6UOikJMxmz71u4pHInOFq5Qimf/8qwLK+YsFyyjfOFU75AtLGbTb3wrAUHSHycy77FfeLSQ4tar
wYZwJwzgXgPsNEJJU0orrwVjYQ+hgKw1KyZFMAycvaXtV0yaZy6L8kdDfP4TvPxU65/O72rQBaK0
5y3Vj+U2PESDLIxtVZ1HhcBwNTs+GJK5yNFoJh+s/dHlf49hgCtGCubym60p5g3sFH0r/xbU0X80
+wnGW2rPPeizHT4+UsII8KPYa9TqnvjL8MXgeiv/vGJh3h+Dc86YBCv2sCsqWSdNzDhhvMJOGxlu
bAsXkJ5ldY7+JdXPH2WKS/YZA+0C0vIvQmRI3ZYlsnMaVHSMasVvbws3Iw1oDFAVFjb/wdqGvukZ
9ZsdP4F90fW5v6BYxni+R/THW3cJhoDO/Js3LZj319OV9Bx+2ZGB6XHkFiLzDfJKf2JlknEO/ZzA
oFmrXRRsL5iYGe7Oed7eKO2dprrt+rFrsVJiStFMGr/Zctm4MBwZdEdr2o2mWiM3ro0nrUM1I1g4
LzaD+XsQ6WnmQ7sfvJPQ9jiloCXEWzu/wSsopyDIdt4w1ZLzTwiz7h2UUT0YWWiX3b59tE9Th4ez
XgOr61PIa7d8tKKaDmEDr5DkyWYKkZb/lQQ1jsqEvWyI63r8aDaXpxr8HGIoG1HdMw+tLBai8Tmv
mvgWBMcT3BnaJj+YcU3qivO3y0X3drSCi0LOI5ppdt5jZ9kDKXs/WWTdKiAVb2MEEZAJ5FUO3Syb
L5Coh2y5sX73xq48j7CSvKglWD6Lfo3K1mNkczJWrt8JlRFwrpPQIZfHZAqRsL+Vb6qnfHI0C5SG
dLumzYyKsDRWWBFkvejaugRBlE0jAyNr/cmvYrrU71BffxY7rOlY5i1UlFEnhizuP3KIv6ltz+i0
vP5ShGw9mj1hUfc8FI1ku6MIm9mvls4KR9WmO+91xN8hs4tDKhsXRF8TnHE21Z54mXchkjo2Xq+M
US2BzP5s9qObAAYPEjrbEfEm1m6bvg/NymZn7mOiGMwS9EfaYmaznzODyf9RIKlBC4TGTgYhwk7N
dEN+ye0pwLdR/T2ATgDhxXOWSNPzBAoVZP5kl7p+WbREYiZYZbGoI3QwQ8F8aglA0/TO4aD1lJCH
QF8wzc5+7AjvW0MGd5dtWlO5lJkAbPD+oz3cyPC4rvnV/Hl1TA3nMNY/T8NHL0eqvVha3ASiHK8i
Ou/UbN8/h+6sXaZz7PyNXQwyvKOgvzBuUU4w+rs+xiEOd71Plo8j9QO4zyeTcv8Rwrt6bUW9IewF
qt6iAW9v3g+wuPTdDLr61dp81YQL5/GkoFHVJMVcpsf+pSzlWMPZl+AhgrOr3aGwiJHNu3FA/3AN
hFvXC4dUgZ+kPkGc2/igXVZGOT+9P28H23NGHJYx6//XCgRkyIBatN2xRpCg+7MHlout3GIGhc+j
C4et6RBSA6+QITFLf3u0cja9roSJgNJ4TrjvzP8tCs4J8hTrIn00rKFVRjo34u4R0s9/D3GaFHOb
lTU1zJxDfCUhKx7Lfv5S048a0o0BF53psWfYI3Nhw3cBDDrXkz0YqMDfKxNj5icvGqtYcPaTn2xv
e7zHO6BGDrQVf3CNKcGGRsRoI+CHCoIiwJEvKSIutblJp3Fqg7wFFs5cABo/8hKueS0w+T3UvaoM
YetJkfqb0EtXAZ8lEVPPh4iW62TTxTb2p4jjwAytQC62nPRHYig+IBFpZWlYmCtWGlw7pW4l7qm9
qXfNi3s0pD9PfzpM+4yKYTKXkGfb8g18O/VcLLg8IkzqwFSTnZpFGqZsiMy9axBJblKupkc4l3b9
O//x8sD/lfe9ivUdsuI5L+HiKRvBPhNUe8QExxjb/dgYaTWNVPfRkrjAxQqQMmCqvvhNJA5Dx05M
DYUrEbn+zfijliudNDe9hFsMCpJapVzLFcvB6LyEh/+YufI338j9B87DPgE9UHTquB2SmDJjP03H
3F+zzW0AGurqsXNdquSnbjfIskZX3mHqs3xDgdN80OVNdOlKTpBAXroexosiYvhGiQoJnk5rfCqY
jdRvZcYzawZ6fHt8AYcavBzIJl2D8eBq4Lche4xuqFYVXeqj94d1CM8YyPQQTWSGj4VksV/XAvug
jZ2nUfjUKnfgDInj0VSdj2zjjYYiLHHL8tgKNbIZsSuNMpMKogccfEMCM3jhm8MWo6bcOHVq1Qbn
4yu5DuP7VaIxrZdLTFXZcTuO8rxeTpV4OzpxF3+qiLE6DipO1JHyS8xXEEdO2Iax4ADAkaI21CW8
f8WyV4qeRdPizK7i68MdhXLCJluFdLkDpGd8IW6zQePkZtGuJP12aqW7mM5pay0f9wpI2LUxs8LZ
JbmA1QYw5L09ZiyVZhS+4NNcndzzdrzwM5tSizeeQZr2O11HjIKq5VLMeSNoostWdzRifHSxs5I9
BgCIlQCM4Sq2haAMaSCQUzT0QIynWIBO1vKitP6PtVmTCp62lfGq0JQZjjj7DeI/RLGqURXRMz+F
q29OhBSO4rRF595YpULN2jiSsL10nSU+zLwl5a/w0CTbExzqVTakjiakO2wQcrfXoiFVMb3CR6Lu
i0qXdhAjxsSlIKft0AmqE/2lEFj9n+c1zYt38BbpIeKF5AGOEB0n0CljTl0EBzBlAdVxsYnfkwQC
bsNmPXeenV2j4WoiPR6urx8OGzsKnwAzr5iAMma93+L1Ce1Ma783WPK0ZCeJdcIc0MXIA+LkPxKD
jbShi+5PzbY1KtV8YExZH5WXXXHkId9LWY4vRZtV7OVxTiFTEJHFApXatY+r1FsVXB+MiEyRxPPr
DFSlBPba0NxZxUJXw7EaTKzeHyBG7RICvsSZb53rXTX5BkqPhJ42bvwc9e4YrAsEel/cqvCGhpQ7
DegOhS+r0eEMeHRYM8bmgxvbHceNOw8/ZTopNMYoXs3pzJXGKMce63A/X6whnX2ajcWvsiM9UDhT
gR6oOA/4lhf2nn+laJa7FsInOsPwzap6g9ofdviTMhLnWYz+LoDlPFb11Ez7gKMlo278OFFB1nkl
tA5tgygfU849BfHC3kDqKrJOX+c0vd1glsMd8I0P2FbtigMa4TDywMuyf/J5Pfsbb0Z0d0e/srHi
rJuRzGgZik6cfo4nwoCLGYSfSkH5fgm7dqV0V2m+jdbWkBGqV0TgNBJH8XAr/rt1E0o+4ecbias9
dkSqhEvw2Z7mQxtDhjkp0CkM20xDSjyP0A1dh6zU4Maz6kRQuaPQafRDlXnHN6llFz9nXkRLW8Kr
rQRgi4/pfZygVZKALoFK4ImkGw1bIJTylBZav5w3g8tBN9QZ2dQMrt8BeZV5sP3/JLJI0iuLtaxs
SE/WdrIm6zDsuMdQgSlnyz5L6RTnO8na/XBD7/Crt3Yx4DIcXd6HZPZJJEgOgc5rMpF7pdLmxau2
Ln/WeZUCMZnwFpH4b412+f9HY3RZuX7VPYRIxiqsRWNS9LN/TUhthSTdcYu5+IIvoLAYvh57slRY
NPX3EQFYEMSOLWaGqOx46+QdyFUx7rg991OAzZajYqhZD2xG+adMuGkKg7P6Pdf+9J6hVfZPqFc/
zwxnZpJYZUkbFAVB94RSAXJOgLVR5VDCj3uz6dVYF+o3whVPKYAonYQa67a+OKzMJjGCAjN26cf5
hXdR7/Kd4aq6I6phhwKLA7gT1H4PUF96WCW7XrX9ZLzWRGxJGzE7W8EGO6zr6MLaehgH5cxTqYxD
S51ZsHnQURyDMLVSN65hrHL72WKHuGMbpPutk3476EKLrCOzXsfmqYE0LGqH8iaDBj/T8cQM3Nvv
ogCZG2vYnPzWihd79w3pcSbetknpBFSPxHKp7Q+Lq+mhaSM7EtsM8OW6HGRilPyW3/GSYuBBoCb3
7Uz7UM9DBo1gCWKH27S+kcRIOg0v7Fd2HuU++85rtlwdnPlARNPd7EI0HaQGzFMi9zWLfkSLUiqf
B+86Ua7nXl3ITvOXD6E99rVwmoNQbI4CUe3qFuf5cJ4aOJVkl9dxdMQv8CPoLYsjFMijCeHDRGke
mjlewCYDur+IyGOMOX7zCPhMsyzYq8w/AHEsztbsNkINWOBffEUgif06EndoSgJaA3Ci3+7b7BZ3
Xi1AlSQNQDJazDwnv3a0ounmgFPp7if4etGFDdDP2IPbVj2htD8oNdi1pjE4I/gaIVGNFDyYFFS/
Jn2dgW49dzlKwYgm067TzYaqeSUCsS+iNuPNeeJJ8ay7EOurVl4dvBqF1hJLXs2OZmwfenPzzwLS
9NYcn62i6MSN4zbU8Ve2dZeZ+IzAzL6qAX01VZjR9D8Q32RtZIrqoiIYf0UMYKyQP/RpZ9+PzngH
ijENoqL7/JL2L/Q8J7HrkYuoIHJgcdUmfn4goqnbyL7Q/5JaEwk/BqfUpCDKd6k0p4oRmwRgXuxh
gMtyi8pWZQ1Zz2301as64prHPjQoXhrEFpuBFVH7bd/nEQsnF8TnqRnX25OV1nW28CyK+XujALQw
rGwTKy0kbvnuu0/sSTuyG+6n7n35Ora3kWeKUrZjTGNmwmvS4j450q//E4K5L8ASxmRwroFhjBnF
kcsO3hQpzVp/g+SBoG/pKMtOeNcB9fyKpA2dEQEj61jeU3uiwjSNmwD+xhM89gJ/m+MIsl73BUzg
8yOXJSEqIvNVUO2LRbBBrhUrW3NGfxZ0xh65GypVS4Esj9ztuvQkW+CAIVtCgHNIuowJTSMVR77O
CNPyIOEfmy1tbIBz+l/1XQf8S1th1CIGScylUy4uTmKpdajV4fGtMWae+i2KoafXGM3S0gvli1m/
sl3VJqqU0UrcxVxASsDhdkbczLSb6TnGz9rUi7hSqFbAol9issOm2au+FN2IdBpqjsTF0JxA9p/s
mJOR6L/M1FGES1Nbaxvd7Wr4nQWU+OG0+ExNFJwDT63A49HNl8IzFViEJ4qTuw/FjPURgqaWSsl5
LFQtdnftqsr1WoD5Jnv+uZWVdfHJjjhwz2aBGJAS94t9fn/N6sfI2rTMEqNax9jtH1ZPI0o8mKzd
6rG7mDCCiPi0yKdtCQsnRyVKJdJnpf96PZwB+4pTMNjbWor6wJjmnpM4a99MW4HqXVG+ATDgsW2K
qeTTLKywhsRhuuTWLW0TW2iFfrfjKQIld5bxYSI/BSnTf7ekPQhBCneYgkMuT9Xfl2n3oe1GSFD9
nws0Z8piYp+TDktc+jwG4GLOxb2fGqCR7fGDYruqjHS2I+AUJ29SeDZNZ7kABO41LxcGqX+BBpyB
3UHg/rTjxxty7xjuDW2badAvWPvF14pETJHl7mU3FVH1wRiIJWVz/Rf8gALdh8v7Y17Uo33Q0OVw
XaU+j6XxRWKhh6Qc4buMpB4TcRu3NWp8X2JxdsM/RM/MGznEb3HOiLGsDYTUrcO9ZlLQedcsWsHP
IRUS9ILHlvZNQj5+9jPMxLdRx22F73ceZqBZQmo2EwsUaKdWrUBrdMSGwbO++Y89Z6pY/2YoTnX1
smuwD2ShSI/oa28FnA/v+CsJNWuSen9pBELPY1Y+i2dmeIcnQXb/vBtnvLdtV8kLoFDNvjUwbvBR
g4D5LGlGMBk3eK+THsbEe4n1+gyInubBULPwnYHW15EKpoN5C5otlJ0DQ0lVZxm8mbGSnbaqeUfu
z/mbdd3fpkaNW2S1LkuJZ4rOqbjoJ8XuBQDLyL8IvYQikPfHifjjwOo/kP8pKo5hFQwnw2Und493
ohQHUFm7Xi+XBgK6qZ3EPInphsdKIxoBgKQfG5UVPH3WdWeDEzs7vBu6/q3P7pJuhYSRwa8NEVhU
ptDa0O8goeJg8ogNc+Pgc0hgkBWGR3OLKFlIjhXAOW25U/htOpVr/mnCL9Cj333QJhdybl1YD1bN
zMqJk9M+8rxXZ8QYCnomS+1B1vkiBM7RveC+5feBxQ1ototFd5PT1iQ/wMztqEmjcKj/PTNTSoFl
5G4Yq6Psr5oz6CyK2LHlfbkC3G4BRgMQhW3MXD4tr6xKc0vBrla81dcaviU7ipNWikW55Gj6twRw
+Fp3xhyKHn61yCcQlwdssxK1MlwKVNQrr3y44BrKW1PpQJb0BD0aY0rsKQ+ZA4rgW+uJOGpQfwwu
y7taahwRL8F/48HvmTpMuEJ32T38EtzlMWaIDF2AXUcML73Y9EyvC9vDHes9g1ti1EqhsA3MwEiO
wepfBx0uPhlXpZm8ZfoKMJe9qZClTje1KwEJFs5ubikAspdROhW3I7WmfqYaOeVLa3ZqbyM1k7ev
IpQm65MTCkaE5NXVtcJPkBIu/CAK4yOICJJbTvTEmOFBRM7FBtu1o+40yXvWnxSpmkN8J5D89kuj
/9snIz2B4UIFQPzX/7d1AeQejw/ezHvAtCy0QW4cJCZw7je3QtvRSWv+vhdMRBz9yQtWtrTEwSlD
ZlRzVW6SpPGYCA0ECZrH8WxIEXusoyk2AVNm1MInETp1ERWBVHNfXtWawg8LvqfaWerpVu4k7ip5
OwrjQGDPORQkNCLQ4Ovyd55e2ITnZOa3Q/bcl3TgIXBQeVKfZFm7zcC/q3bewL99Yt6yZSw4KvDG
oQkQfMckiXcwV69+bz4RhfwZEqmxlpdkU8CCoKgaqy6wzUpreorS/jd/UkUuD8tDS6rWBSz5cREH
z645/pGSUPxLtuAMVuA7DMxcqvy6rHaraoSTysj3zrsge2rh6fpQq5kVJrLto86jpSGNyk7VwHzy
hNx/4IzyZRxxC6PtRSmGZ4cB1AWr0Mik0BMA8pmm8WlUiBAwgGcc52PN7KY1SACseS2HTpp/325R
c+Kc0wG5euGDxAeKs1nOSkAQF7pO5oAJhwjcnDkCwquq5E3/9Uxui44HVBlINhryAorBleYum85A
d0RS0RS2PMidInYsUIpYNn+Wud1N5azMD40Co4LABd9Inwdii5q49itehFSKWBA5dgZPGQj4RqpS
osssOLEf7jCbmJUV7QxjOt2qz42EDNrrTK8nzjxIgDYuom53a5ufnGJKPIcbHK0G2r5M3a3uPDlA
UTBH1FmqCklNh9R4hhlOK+fNCWxtf4niyVtH5OuS7GGuFoGbUfUM6Yw3EscOq1qgZ+SU6GSEHv5h
MEZJb0G2GlTp1zcWC6TnwE3GJY+HvvoNr7vgD2oyL70PeleKH+xDACiRxg7CHo5kgvYdUfRTGdtM
ThvlteYwpVZhCFe/ytPsIEx3JajQCuxTbxSVFXvWsq0qi7hqUqBY8N09tTNHj7mcTTowjy9o5Ssm
U6CzOs4BsqWC/SfKMDg1QT8y0RxLLKXdLjsdLUKfhB9UfwTG3FU7ZFxPiWmCBJp1u0VlGvRCVFGA
djK+S6eoBa7epm5xgyLFIRB6h+B/6c573OkyoOdkxZ6CrM4p79Gg+seItpFl1gSWUcdonrTclye4
V7cL7CMDwx+asXvt0Kt8e+jGt2qG+Ckli7rCrxDC8+o5mpkozoZqVY7ByVI6+zG+9g9ygvsrFPeb
Wm8Sm4HMEZhGDuiaJ79z5krYb6DgFMc71Gul3zGUmoZN3HHmQwWZFnBaSAZCKnu4ltF/U4zhulUW
ti5CyZmb8z2z8B62mLbBBCWhA8+pns+kZFqdny+jBdy+8nXXa3Gx/YZzidJyMastlevRhlUFHHJF
ZOXFNL3tvx1nGU+ReQmS5ROVUz7HDzXCApRB5KL1SKwkCbpxzK9eJs4DIQm2Gugxs4F1hNhMdobO
EAb4hlAJBaI0gLvWWQAx7JkLNpNtfh9C4P4QVlCa3tkYWCdmzmT1XUEUKICnzSGaptN+b5QJNuzv
1QR+O3nE2qAQCVziSkanC5DIy8nnPqtI1R9Z17k4bBjJRkCxkVUyKKg16jEYgqwHtLH5RdZHLiW3
G8NTbogAnShOeSYMotg3TA7k4Led0yJ+e407ZWGdm1KzX9vujDgvChsTJYDyE3ojUELUi6u+zdeJ
M9Vc0OACOCQbvSQw9mLym52LWbIA5i+2NrE1OiFr+3pUfFjTI85JvIApFrZwxHMTrPef8DvPzw80
0SXcKx4DzKid1XzEaxKzm71et94akQSyb6vmNUhbq6Iqr6J9RAHTAKp7v+ZMzegRMyzd4SV/pTw7
wRmYiLRIEPZCxeyfkqmPB4AOxQ8jQd5LMvmQmNKa3pi/hXLGCsvetJ4mPMN2jtqxnR0S+Cfn15Gn
hc8NWTdOfF10PCfxLk86GX8EyOvjUJPmaN3bwaoCUSQv7/EdRZoVZBZNAQHaKb20VAjtDfysZxFT
z4COpCZhMGKhxc0seAIN2xTvmPDkc+9M5+Sd8lawfjS4fsP1dwOz36nMIhsSEYYXOFmTOcjUTOME
aND2oDed7EhcQ+IV5CdfwFP5YDCXu6IGvd1zfdUSLr856p9KRYtI9S1mSzSjsCD9rMyn/92+DHc1
YExrm6Oec4XxIxqOtXLlL6ROaHz9F0ZiFWjz5cYnMnp0dVS5Q1bnK2Uu246aYZEiWIlhWHi5akgz
Sr42UK96DfMguHIDepYkDEab2GlmWgDBSmv0wzvl+pmHTPcgOOsxsgNkSZzke8Rc2Py9lJ23uekA
eZfcsrBRo5STbRrWRdiHxNELtv63umNgD+LkzHunraFWwe2rklAWuXH2kbAUu/gwuWsrp4JGfRgM
SeIKHm4GyIl0HdGxdqpik/qXOKVBpnYlmZJgSGo20tJICozS6fScLXgDlqJJ5vosAaRPcho+Yl5Z
le6BWmqKeCQD+8r66uyV7iJDNhLtNa5TdMK63qxqS6Zw9ITuCt534SJkie2Fg+LsvRWRPiBbUmoX
qoJFhRHB2Q5jMdzE9X7xCf1n4zlZhtA/pE4OkgscFVNRNah2JTbndHj0qjRzU38n00Z1N/SgAJ7z
QtiHxh/GLBpMv7rHZK/bU35sINq5ZESOEUy2BA0aMhjVURN6jNHazkuBG16I1dvz0t03rpL+VOvd
pA1c2U6OGONoy/os4KOYdMiTnE0htFMB/xlludM3UTU1UkrbhN0J0vUALAiUpuAfBQcZqE/fKgBZ
ue9ue6GLXKvH8K+jI24QOV4gc32eVy8sHArTGb3OkoaB/Jm1PoRyj3cKUvlpYRKEbeYR6LMkCGpg
Ma7Sus7OJP4hO1eu78AvLED/yWXFNNjIXm1+JeXbHwAZCxRcZk8MxXhz2Bqx5qN3bNBQR8VeHjSv
4Kzryx7Sv+R3vvpVZQZhXFX6A+jKEGB10Q08EpEOj8PhdJ86EGe3JN8k9R2KRiI3D4hi93rAksEe
yuxZqCEuf0JkMSIkVOIs3wKEZi4gkCMnbmDNMLsQLG+gAtR1Dxm5IQwVJWhvlTzGX0B1iJnBQ+Ls
3CXliEIWtxm3DmcEEJUdhu5Eau+HmHceV4K1TB2jTUw9P//Nw9OeagBQIAQDhp8/doxOou7IpLK0
bE2Veel/1LNwq3meUs5y4qSc2tw1WvTjOkYZJnQLyNQiCqtmSk1AZGs6x9ElfLPOB7bA+FeHnTE6
MfRZ9nsMRlDlc6cWq6mG7bkSwNy/WNzuuAZ1rAzJJx8ZEgau9xdnR23EcT8SGK7jOxHtI22jWvoM
72nNNtRiHT4uQwk19Tz3mPnhY6Q27cyGT8at+AsYF6tt2rA2lhcw4w/EB7ISnveJOqTBaUfSb1O4
W72MHlg8qHytE8WpoJjih3SQMZW2DgTCPuuPU9StyYezeVk4uVMOJEiuGWk9xVrboMkAgrDmYkSm
xjaGKqxbaqqyuQhJ3BUmjl9Wn4q3FPZNFRSgA1x0jKNr0YLD8orXfs+58FKgCIwsiHYNpr2vwWIP
jfIwpLmyGvfPCoGoZlZf6sgtTYmNxtJVb0pcr1NFNCTuWJWLIAbej27wRj8LsklJj/b1nP/0y1oa
FiVpg+38+1feFrNu3ucyVWOj/a17Bk3oBeC05zNRD4sgoU7KvLQWFJ+zJQbgZR0KQFwZgk2o712k
eVXzcvUMFqBTN76Va7zKfJZY8Ba7O8UaBQbop+EZWZOfXy4M9XQ47QeCx0E4yn6NYuvlmaNvFOWB
ye5gDTuiFZF29QFyM0gD1zxjT1KrEwuorvo2hEFP0JlZpq4RInGewJeazuS2sv0l2B3XLe9sjG62
xK7UmcUw8SFmAT5a+0OPnButvj7dTOhRjRdH8Z7JQrRXcvnKsBj/rLES0JM5w8JVOc4m/FBHAZjB
Ibaj3gJQ/llmGRLVyCrtqX8Mk783l9IAbhFkitWe5nJFfa+amDj5SKcGE+uLy48d5ii9kmE54jFV
ptcaf3f+5Ca77w8QjVABH2MY4NRqWgHKoBItfHvmeYYZfMG66PYXYpNNk+hvM10gJ5o2FSy5wuhB
9Kn+uyBrFqkmcr2jhM8denSuzWG1IU3ziDVEtbebKGSvpl65vqTOb/15sG7if0iCxZ+OsssKAWp8
oW5FgcCCQ9yAIOmSGrisyVrdsoeC1+fO3i/899Tv7NkOnamxfjZcdqLkbEBKiUmRU69raUDe8GH5
yu+hZld6NTjWN0XTXKYWwY0cEoaEzB87YwYO/ipHMhzhrOqSPIHQLt3Omz6t8lAqPjxFJBBOqItd
QSQPG5PAd/B3WQtf59hoJGpci8HwVM69jVijAlkaMP+Ms4j7S8EKQT19J1hdZdlZdJhTYUgL8xbI
Tc43t1I2yoL0S8nChmobGYa10lN/khZqnLyl99ao2vLMfW6/NsXCIrrCmfIv5Z8WBQzDp4HK6Yz6
YY9yn1QOeUR8igEby1/9YVEw5eV9nlbDu/OjIIGY42WiPiCSr3ZMfVnzej6C4RLMkt4yYsdklNG4
pfa+W7X3RAFRRzKbFP5hjDVtyWassBImtW5J15e0D7OLog3iqs9DZOgiwJ+icV8fgDQVOobiWb2Y
LMiINb3laUFg23E2qvJZr2/BtkXhQujULxxpct1gfXu2s+3FIx5XeXpjWdCoznOzYGY3OzAqsoHB
O2TmT/LkXaI2saAFj9lFwrcImcSS8YAJwxxK2dJ5UlewCktTw4APSmy4nRE3B3yKx9gSKr5ZrWn3
B9KlC0PncCAGGzQW4sSJoWy33Up2WvEMQFL/iBT9wwQGe4ETkGfT24h1JLtpMg6dXLoKHnbrQI22
HfMgMovbxJyZKhtY5DEwsjqaAHTenNGk5PI8OosiPn2qUxEzsb5UoRLjfrn0ZneYmeC0LccPNdzy
yLS8HsVy7OmzFYgeIVsMryNILzBY+y1OT9Czda9hWhTrQlPSk4sB85sxsSASlVaUGr3WCSuzVCQc
9cbGZA9jIEu2e9Vn25llJId/1XBoqBV65AeLjqJ7+F7Q/JO1wjfVN1M7ArAPpj+Hwaah9T0Zjxy5
0/OczyLqx6Wulg7Kr6BJ3mHXxoTMAgjzp3HaR8Ib1YTQZBt8bnz+PUWDhg2pDIorFaMbzZPUd+Bs
RmgauhMA0O1lDLY7g5tj2KHvv8xLpEmQjdPP0oTsDnaLFJC+zxIqE4w50B6sDl2xooBPTkIKp0Lg
VkBRtRScB71yACUjMm3UoEuqziiSxNy8yEraIb2YxJFiwRgA7VL2q3AvY4daBo9dQiV8QeHmri3F
DYpPA1QRQP9J/Trrove4DNIYwH4OnvMEME7SFtomgXxyOPmqf5iMwDfVt45MLezEypB3DNjyPmsr
o4W0Xsg8RQjVZGLaiZ1x+KSjyTDP7+K1yZxJwZYEYsSDfEKDI3nMF9NxUU+iT+z1jCvvZZUPdJEA
MoxwSrcD8t/8PW1WsO+U4lhYd60yHeD0SRzotqhbDJ/J+S905UweOso9LcaDUjumPSt6xUS9G/kw
aSmXTA6Hy7Cf0M75ZzbL0Fj5gL9VBMrheJfYKm7PY4jfQND4FUnILr+VkBVgiYMedLtiq0F7J3Lm
cyzt74q9ugYJ7yo8cLdH6khpjJF6bxEcHfDjtCCj8Y7PAo3AcHSE2TozxIJe9VhU07WAyAmauMnM
vOA7eWAlQBLPYHEmmBYVhfS6WU7hraRUF2Vdn3ctiMAprid/8UwlzT8KNmVWFs9KtxLJpn0KBqvT
syJq58GzI/6lLQlXsuW6IexMQY9shGK+zzqU77EXxG20eg0+0m8ACMws63JOek7sEt3UumCgc9BZ
X12DuaggT/xf0VO3i0tKESaNy5gpOUQdPkcsfq75wRPIJyiOSfYVUHgXX3FWDTyVG22k1bNTXTkW
pAXL+6BLKbMKrU/H0Y0haav/DfFkevOq94Hu4R6mImWtkg3AjvY/jr+andtUTbfRSk1L1P/RslUh
WoBa+WC1O7uQ8lj6wDamKNC2cs2BjC/z9LLCQtMnifejENKdKSTETmxU+sz7sq5KKshb2HXJIXov
8uaNOH2rhEWFOJy6tM+BnzaxwGAokq2jE6WB5R3JlnhRzZLfriRlweLM30rJclZpfoM/PKJ38q3m
XJskaiEM1qW2PfAoOmu4y98kivFD9uYS1HktkW6NZ+CSAb4jCzJtLGC3JKTa/C1I7RlUDUVcbNjR
nlF3ooqgJxLH5WBkZS/IIBmYclz89tQpIQ4YXC50aBL1RXj/1UKlw1oOIfxh8909hLfFZNtnGhV1
DUvUTr0o9Gn6RlDxSJFcRR+ELIxqq1e42DwzyOAJltsoReUx1tX+M446ANW7Q1iHM3rJe4MdKHUf
coanmDmCPd533eKnxBrcXTte8WszNXVpRoGIoUgRbhklVIO9DlIKs2fCrMX53Gpv6cLhTNZqaB5U
dOWpsP/N36YXtYOTJCR66QdZQR4g7bjPm/VsnIiXPI4HJ+oj/rR9KmTZBINotWhMei5hZnq+iYjo
WKMWo+HytINtLDWxiMfg4G22Yhx4YPVYqsRsAr50Uoj19RuFYarJFttTKp1DfQbYF3BOOezKgVZd
y5hRu7umOILqLN4J1y3nvwpA2N09IJLMrcqIps4szkqUkUOz0CtiYMRjj+ga2RWLvpfQ87pHlHbx
V0hgfs0lBT7gM4xmljw5sqzXnjgX99TwIGGtegNav/AGKNSIgI/leAssNkraGBKGoP6Af0mNVKAp
7DEiF2YmnSfkz5QIn9/yryYUZEDkJSFzb6F4OzasWTxBd2OUt4gCXG2BJzqgdygtplrdfPqcEZgP
7l5RL1t+MWj/R2hlZ+TvWXPiIwsEwdGuo38SJG4sqwkeHQ2YUnHftm/G5sBTDALW7CwDHCM9cfmu
o/yuWCDZkUYN7ZfmZ2lbUxEpuvectBjBHLc59i9NZJXJ5ulE/EOdoE6dW9hvEuGPt4S5lFhq8dR7
9SHT03UMFQ+0u9t5CcZNjpAxCzv9AUSxj5oOFWyGUqlGQ3qLk8lC05NxJavncU1A13CBU+CTcfbu
EwCSzYI3IYfE0qrXclQBBGA7GfGX9yjn6spPp716SKoRElFtDBQl+xiNwL018GzizaU1YQ4/AVAL
tLXg4fxDt9DnznVz70i+jCyiSBkNDgJeZePb9+VXvXGT8J2ice/7XyYAoXh4YWkpKpLcYo1RSAOO
aETirSzdD1pIvXtQ4kUAmFU0XwZnx4u/54LLYf7Uu5GhDP+HTrRA+d2mwgi86cPoyrz1mWD8bbYc
APoV1mCuX+EQxJHyGwH6FMvBQ5AFw5g4xkvR4H4FC6yAhFIubH6C35cJzQPT8o7RvgZLLMUuywY5
CVv3VaPLlPizukqo7J7Wvri5lsD+d14Zgu4B6jg7AysLAzxkgATSKzL0O9yABESlt0+Ev1Sj56Sp
dzMj8vw0RiHmIXiS672m1y6p3GljN+6FmH39S0X4yzhDEQ9wn4jyMWos6DOGzQmtjmlxnTkjV4aZ
Egi4mAFBuxhYwfoop+/o6oYZOxcipMpIGFWrP9eMIZREP+um0XpLVGEMBiVPaKQ/A/zXQMcCRKPy
wRvfamX/cn8pxKPorrzMynPyTbw71fQhKkfRhFylJJNPuR7HM3waEWS6t0/waMrYbO1JmefHMxat
ExUhCE3HjnhblmDLQmSA6DZjD7GcxEaIYUJaa5kt5QKNRDnPLBvsUAfUxLP/7ITBXY8TYyXPVyNH
dBijCj4XWY+1al44+Nb+5FtVll2R69CMljun4fNSA2J9fD/hnBuEd7/qG921JzK7nKYqoTXvMIKw
OJWi5/TpVNh12HeBA65ufKAY844PcZ3oG5rXMc0gJCll1WgAwxM2qrtYC/LRmY7/gCpEeZ570ShJ
TirqWHIeFY2a3qql5DlCRmUE1FdEsq1xjE0dDgMKtj4as6I5FQ9wx3jiz05fOxPBQmbSJg/FRCCC
cHD7kjFdirCD9W9PaokJey0aw74PCNqm5zogFMvtN1bd/cLWx8LVcnSUP5ctoKApvUs3uowzmsG+
N1Dh9c0SNT9L3CKeFhVsbCtZgypKIKZTCMJ8obYijObGAnSX9OZtwsJZujwfHOdeBN4chADMzLgY
MmrKrXhVXHp0z8wteeQDWQLybX4w1SB4r9t58uWhbCEi7srmH33O0ew9ZtMtXBmEaxkyTR0sFvig
L23RqdhZnQrVxKvQozsLAHfm9BHOFHL9rOIwUeOscJrHxlHWheHQn0CcHbWosg5o4kgAwYXGiBZK
FCrHBhs9J+5IPheQs9n1ivMTtApZqZ0UF2FcHMliSa1qRs8xvExGT4j1FIxXebO3/xiNKzVxw9YU
eVi03F/v26gM6y4YRlF8X4aHYwBgcNZORzw4QnNmjMvcW//Iv1VeD5k2CGoa5RjCp32Ggd/H+oSH
tdOYlVVX4YoWEPThnFBFg9BmZoMjWAK24RWKPzgtrMHaK1l7xm/8AfVAyBzOg3JfrQT+IGNF4deP
+YJ1KlG0lIhBJQbYY0pLeL1SKizup6rnU4kk87h8j3WXlVwEUCc1A6GIgV+PrnZAZXfH4oJA2Gkj
qzwxmUCuPHkePyp5ErJiaOuNjyEruAT/gR/q8eN8wYLYhkY9RUWPW0EgetW9Eqiksiho/rEXOndM
/wP0TfvTsRwOwWVeMuMSbi0fhEbuccO8QiWABTmyLMfkUmtMAlZJPO0UrYTP1F43kUE/tNYOeZR5
DMq86Oy7UjvdT1lRWU00Esd8VPawQby5I+Uf5MDkKldYlNYlmn1nZpx4JkUiGOs9+6Zp2UYF14Y/
f8bdLLSKiwsw2bs5852hhL1IvmlA5jO9P9R+0ysZTWD+WOvgSIeh4qTh/QQiydgPJeDABlNi8ZPa
pdCd92SSQCRFsyFwVDuNbNIAyJzdK8mpWs8R9qbqMK8zk7N9Kt2lY7/ErlDLu4FOusIisiZhuJ1F
n8IsnGS3Grkr4o+3VIH1zsfpbX4g/S2W8prJE+kmQis/3QrVpj44If/4/tzG3SmPXgNRq1KgLUym
8PxKJNr46tL0ng/B7iZHwOndh/qPA5q1uF4kDRHJQbs6eB20jvYGvQAQxWeJjFJnUv8ktwJfWSbw
Dmp0Ko/MCFGbvVUszX7KIS5kK+V2k/bta9LgG3cWTSWkHFcsEcW/mh9gsTOO4ogmCRa7x8BfJv/Q
40khNO919109jMMmnln6ibeeAEBCNfkL3l8eQcjQKf1+cRUcjLhFCzfD3J+VErQ1lZvuKT5ZkL4y
yLLJ60OGBx2cS6mOa87x0A6JGq7TnKLukl5wb450JQA2MoTtpU06J/SKClueHVwXU4A97wN0AN2u
6BDcTBT8TKj7RutmZm1sXqh/d4+GqPaNfZ0KntCXD5RgaGNdv9+1JQr73oXY8AREbYfgaDfyu6VP
YfxBxo9DiJgMoBB5QRHHqdQZFwcNl77XW6WV0BrpoCjUDcSq1PtRg4PfUqDBU+8fmu3nUGkCHy9m
k9oYYik+R1yY74kCfwB5JBJ0Kgrf5/eUZXQBz3apUSCl50FqsxXKzKvx/wvGoo3gbL7CBwCRoFAj
30Ag/xxxNhqXUG7YKYSs09YASy3v6yzWhHPtnScZZgng1QZz6Qe3Itgk4ILkDzP6+G/FB5G9JmHH
SRKdimlvTy3zWEBU032ln0+mrfoZ792eHEjJeIqNkniHEfqpmPJx4jTqv/Mt3br/3HIkUKjrBNuz
C5aqhkTO3WT1FTMNrB9M4nQn2LTAs8cgkaEdrfqb+21DjyrPok5Vk/OMR3Z8xBHLdLNbRrHdHidX
3Ns5Ic4qx5dejUw89IqltUXgcrjC04CH1kXaDmi65EGCtxXqsXugraUq/fgTtWeqEGGuWSghKNKE
Wt+Rn2sEsjZSxkPz/+fNxRCVRM8iSUiIUzrvMTR0Tzt8srJ/fM4PyoN80MQ+C7lEDVpbZMzI6Jk8
NZxqHtnZRAPnpXUPkXaCiK/N4L0M5NBGjIhnlR70MNcOvLd0sWh48WzDcNFT4pMNajpv9VMmZG7y
YizriHYpxp1+UKtzw4HiWCwt4vbxbpGZR4rs/z1IMtg7OaF230izW6R5JCJDixELwpIRGK9QfBYb
gLz7HingHEuHcjahe7wLj8vS2THJByLVKHkKpdI/yzqzpwvPRTA+PsAlWBIaQHK3KKljMDiz/VLR
M+ORs8jvFz4hYxmJ7EA7ORkFF8bs1+UdH21wl/qwhYhLkLmMcGwDmd/qh6Xj8CSdRVd7ghCNKSPB
woqOTfq7EHJkbEUXOypnsWYN2rXGXY3isiuEfZfI3OeAr6pRrjiIVJVWbGIP0BEMCpxZnDdQ3784
Vfe4eYwhPd3ul2e6i1DDawF2J5MaoSIWKGPIoVaj33bDGRXVYc9f9ahxXsJ/s/QL1hTYp9z+Aw3J
cTi/8r0N+k08GT5rbtVtFf86BkseOD6APRh2pja/v1mNHFo5u3hNFyxHPOmZFVK3JrbTLlL1L7H0
ev2FlEyxjeydeHw4ZUWGzF1gfAbOj68aZJt4V9+BPXqe+iT6QggNk0im9i+sFdjX3ic2o6vMMRF+
SdtTxUuXUtzrQbXSGJi6Z43XhFgsHV1PZTbVbii6zJ79ZnpVua9WiErTtOXA7klwPVdtYnwZyqKx
R0b4TuuaatCOvs4ODZtlUt4dyu2XQjJBPg1WIUeSRt2VbAzCf9yw3OjMRwDWRAj4sO7mUuki6jXj
WtlatrfWDF1H6LI7cQ5Cvv6aPMr/8OclFYIin0ZCyxX71pkCxKBjShbEYrExy3woZpx6H66T92dq
0/bzgZC5Ax1wd0EXUuanAJyPN8F3e0LX5pHh+XSVVjTtBKGhHHq/7A+3fBfyl1ypr4324lBjC0WA
Zq+IdvNrz8meb6rd2AvVOaNocm/1SIaaHGsUMXsE5bAuS+eG26lk8pmH+ipxoQLyb6ZBpeY/X7lf
Hi9OoEIC17OS8apYS5yB1Xx2jOlLoUTh1IP98zYK1xSTxK2dduQBdcReabl8AuB16/v+mvv+E4ZG
TCaHlp01orz27GCz3EkUE3uOB7g8sEdrzqptjlyQBRtAgI3uMbftXVO0BCX4friAPRWKLQ24lDFX
YNUXAvvBTOrn7CIlJOyPtve3qbnFg19Cyud1pPce4t8HuhNGmRKWht5blRGZw6AqPsyz5dxqvicx
QfScW+MGMgJ/9aJw8EgZ6m4nQUY01gzSHcluYuAKkALoPbv/p1LDH5harc0QmdgZQwoh1Vq8+j+a
pdLRtwcdxfSH1c/0GFDDIYrIpBQBwYqpKictURdWFHlZTIL/JfUuErFowfv5R5kClKu9zy9pl6Ty
cDylebNlzneK4aSxK/WMoG2DDv4E44VIdpdaiv8d/Vlx/PYocyTRqhDEKKL3DoEAQ6Ne00uv52xN
u2axhWF57kNKq0J+dFJ3iD2OVyJ32jziD2cU9ORQzypNPOkRlQcowyO8iZFjx9gzkG/mGL3CX/16
UIc01StPjytDU5YHLMWxx5ttkY3WbbBK4tv1kexoo/O5mGbO6CAI5AAn/hqtIYrtS7i1ehQJufy/
T/U9xBpoSZ5msrK+Z5hyp4lNLTnKRoVUaF+C5D5wKGV511XJFmgHXi5jg6Myfc37cJnCyLQ7HWMP
G3PaXQEUp6YgzOJsxt1GStD1IbGiWQGr/F1uDnkALTIy5lOAROIyk54VVPyauabK3KJM3KiM61/J
FndPruaysVhLROSwdAL8OV67G7rdVl5uBnS2ImqnRfWdme6YJr2oCg7Ea5eIvkZKfY1GDV0yZAGS
7IbchlcSJOtM9CWTj2p2ZH7eOtEnGdX/GfQktgRPfAPWNo9ab6/qHqjwAjEAVtx6vd68TyV2U8s3
yWHe9h2WEhHbrjB0RSHHr4b/NEZhaXwIHTqr4Vu3iWnJ7cddFkoB1BKztTiN7spy0y3AYaIH3cnX
Ti822DbAqAkBxmewE0a5Wl6zXs/1WdLkg8ZGcIGqiEpJvvih3kcJqTUPN73fLFiWFGcezXsDxCM6
dAbwUH4iJgz2kQhHN1I90Nlb9+m2koWywfiUiDbz53UWQhYu2p5uEwG91yZdjQSOm0oYgbNMPZac
Q3SKoRhGP8vmxCY0T/HoQGRoxCvRI9QFPUAdYqt8dpoQwHK9lnHGelurs2IdjLMPU0x0voRQP07E
RoDuiQjCqLvnde71d4viqCiO44V+fatUZFcHkLBLWzzWfBJ6kVeoidpdvGjjP8Iv6WH9XzvFcrIh
MdGGr1a6hD5qDLHHdyAijoduqZOF5t1P0JYZ42eP2Jq9lT1f/xnPeLe2M8ed3w4q/E8YeD3KMSuo
f/wN5ht2K2+D64l9OQEA4xSP8MuREq015qcixT/z+BFVAtK7X68YxE+8aT337BqY0R6Dw/9PH/WV
/Ou8MEv/2a2pJKI2VmWlKfUZomDLDD/2X4sC3xfeSV8vGYCgaeIFWUivznmGYyudfpXPQXxDLaKy
KZxLP1TuR8H/0LJTpnRDDcmYT0Gp0GjsLUP9EtO42GMekMu798Epr9tjXvhBzsJzG+q7i09F6g38
6mn/lLzllmRne+9sNUX0K4uQwgDq0AIflTGH9QGAGw+/2mb6ggRL8/aCZPYFkNE3bpgtTsb0xIEV
KUAMZ64tgUPpHrrflmM6LWHGaGpP+wKNvs8i4qYVpKzNZCvwno/oHYQkBrxk8KCNh/mtRZZfGWuT
kenHhrfTKbPOfNxvrlWzbcaL5ut5n05ugRsrN5Vyiz2o7Lykv35UqhvWejJq6JMgrucAAmHTRmTN
+60D/5xTNyvLH6x7Gh+mD0pzcgMKLaFDIpRgOKzS3vtHFT0rLbDFqxyQfHX/3tXbw3Lc878/Btm1
RgS53QmXAPO8zlBj/XftaoFAUYtMzmvQWvL9d8ycVsYRKtw5g+sJcLYxJ8n3BnERs8evHhfExhuZ
pa6IkfbU5UJyHrGpOLLFCLaj4cShViIJt02DROszl5rhUP5TlPQN3Lk/3WtJVT7n7sxqucoiL4j8
tKJ+OlBqukONqa00CCFukmWcFVOIiRQ2+CYYLYhUo3XymDFOoOEhM28STAlICevhgIQv9270CPJ6
r7nhFTcWGPf7RDnbbUOgZcAPB4gMaaipcR75QJgX0y46cftzqmYsWG0hR0iUevtQr2ZJ1pDwisHq
+/y+ggsrIC2wmOevJXadERzeiGd/Q1apMEgvPpt6X7k82O0YW55ISwqTQ1XhttvEpwaZLeod/ArJ
d21zgLgBmthrOfNO+HAsI4Kfmwa/szqkx3ou5mYI1b4R8BrfDibPnDgJYaegM/s7HRa9u7/C2XVQ
pzWZqoFZWZ8D8f8O9+gJeqZhuYSyjX3OBR/11T2+Zbpb+Vgq5+om0ZTTzMLYRuzfDrFh1kMkwMG7
BBgvIxEfJ0WRP4LF2yaXVJdjdJ4rVlYxm0T2zHPgkz8vbOSCWhiiJ9md0mylmiK1qUyCg/Gz7i+G
CfBsqqPoGE/ARDrLdUFXiinkP/3MjmNX49gCZUYiOxOAQSLwOOyFXFGRbLnnTMv1bzFecqYETWTk
o2snjNhizzEMExlFXtrIK3fXCEaIDzVMD/KIsHxcK02rOSZkPI1tva6XJZXz71mJvL0Ws/8Q3pND
Bogc2/6EvLMWr8FoNi0vLXTfS/adJcHlfUncAc2COg8E+Vcdb1/RjTU5FJdrFqCgT2/UB1buDL72
UXOerXqSKtUlU24JE7wpk/eiNe2rmfmg5/Qd9v2j6EmoNSoYBvnOALszDM8K9JKQRLaT4mk/63I6
MvE9sewnfwHhlnqsiTshT6vVcitWu3JrRIuMo8ih9ApV6y0w71XGtbvkJd3v6BUaaHy+zNiuF0WQ
hABQjhd3LaZXtzLXcLLhYu49xlw63UZ4iLR3IqjMJ0dpH8u8s7F2DclhoIcJIWBcNp5kVZnWYpT1
YNdU0EdYzQHn187FdpAmXV4KOdHrEkQV5a2I+yEeBrD1sqtufr4QHiOrsjC47PhcfHY4zyX5DeiU
CE6ZVv42/ppqXnj2GpnjS2BuVAUbb93Tf8EJhstaZuGLZnyYUDOjB3A0iriV5OKBbiu5Zufh4fDh
TaAKxQHpfONHtONAmCwrPsY2ofzJ4tf5FSDBOLzvhv+vYB1oIH72Bht5sKy6qvZFAV+sAckYTDsM
jbS02wYDgNc3a5oRcENC9DkeM8QKoEKcWVNqeKYMeFzektRnrViT8viplnzk9+rJISQ7u6y6D/WX
EMoDNT0xvZu1THqUlAeo6MV1sbUe6LagtmwkaS2b+5SqeakYz1dNEVXOAWWmT0yni9NhD3Uj7s6U
a3HpM737TI11o1y3H73qg/qi2scQKpS3M74IHb2ZOkjoygF1bqyP/Ii0Oot594QVotATOzCPahU8
o0vkTR96b8QLdvIa5eVhlkpHTlJVZGMm8DBm7Nnn/v/V3m6ury9DQbXCFfDUCy2nbsXFGQC8x2Kb
d01P6Kd6G5PwpKambL3vG8LjAYvceFyL0bP3EaDgvg/tc48M2OBtRbrHLQcbfr3wcvLFL+5kR5eU
Kj8l3kGDJ9gjk3Dhgxr5rjLct0Bk28zfpmEkoIO/ToR6nHo23l6pUX0X7MW8o9O4VoAvPuA60NSf
kaFr3XAx4DWnMSNdyc2DZkCgednCNm+kYhwoBD9WKttkrC3BWqrxufrwvUTwNkFOoaS3uwfNOPdH
lsGwmW2l3tmZvG8jKlSA7xEk1dhgsfQDlZNio6HWSiL+NsT6dcfEpEjWCwh9sgD9HlYxm3715pV7
gcxElQY62zMJVufB/iiyTiIfV3jjCfipCgKKQ5eMedfDTIP26HsonTaa2A0nQYchXuQ6H49HhPCS
MlJCwt0eYWX7V5KcMmUCIwy/Vr7s77n5uf1WA8SM26mcosH/wBfaOIaQoOyoqkh1hMh8Nx+X3k+j
8A8/dXro5CC97TMDLevzJ+E4NnKJ7BGYDbXMB7P1rQPyGKup3+RlGk4he8WSrKhFO77W48zTITPI
8Y8EZnv78yh+GkNH9lUO21WI4zWv1pHZWMzkmmbp8cZ2giLLbyH31gLtA9/+fy6J3S6Tui+2dQrN
Zt0W+AqxMZaJMLs4pToLt6MZbnw6Q+eEcs0qq4EYQEm4HiQYwd9zfV+IikZam6z2sFJ9nFaXS6Uj
rrnpUmrmeK4Gw0RY2tMYBIHdsGntHwN/659aMwuGwvXVZHII4jtyqq6kxXSri+Rj3llW+E6qbMzq
P5WknlkZ1JYJMamHo7KSvtyj6WrK5TTQtDH5BKos5lPHS6fm+9hI9vn9i+NBSDu/3vpCxF6onf3N
GTnKkS+PdOJE4ucIJAzxOM/YHxW41FMnUJMuJQvC3qap1MjqL5f19eubffBJWjQbeVstbu/Z7Rxg
Y6vATr1Nzg47dBsoSlZaeZxbHa7WjaYjQ97EPjv8o8zkftvKX4HJOYY1PhPdvr8nE/9xEriYa6ng
dLja4ePTqNVuYfksHM4WMKQ2W/CknkKlsTvAwHn2pGU/dmqfOAQ+1h3v8g1jWGoTIQMyanHUmQIz
pjz04J8tJXhl95DzOjFKGFB3T8YUNP8zhSaoW3YkiIuDhJpVKJu+1DPzWWHBzTe/WTkVBpFJZabe
AuC6jUWzVFxzwH9kE+pjvQkkcIi4T55n4qQDkLpTQiVpSkYZiN9DGpxSR+6bjBzD1qzUW2q7z06x
HYB4lvIEuPn7VpOJCa5++nvNV7sJplQYLptwpPv8Moh8h2ceC2pXJOpqu3x+b/kCcvKpXJoDXp3i
DgkDV7MUYWTk45vzTbQmKwo8kB+gKV28WUkaeTQOUJDIX+6VIfntIVixrOQnYsuEvDM3z7kcpp/J
LBz0E5Ps16qbRC9q7i4cgWJ2LUrgxjbHeNUQjtNoapiuxHKJgdHDYUsneu94RY0TPWkqOgSOcml1
GRONPs/CBy/x0Gssj8RDVmZYELs8FDXA7dE5ZhlbRI5jFAf+HAb1fWKbiapxIqSbIdtOGajylnW7
1mMIcj1SSTiC+X8AaczD1d6Vv9n9OOWoRiSVExZfQuXo+gOlIvDYXvUVAvR7d7uQ8uWMkD2LG7Jw
Jlg9JVJakN4+9p2krcdc+dL5u4dWLfQSoM4D3WnI6X3y4CZmalOdm3ld7xao/7AvtNUsRdJRfrTo
AhBVm7Gl+4jCLPrQjcvxjsGw6se/f1HAV6JIpP7D1Io7TmXXmdz9h3bFKTvfqQLEl7edkxQUnpI9
160fwhxMiFc0XgIT1oHbfgMGiQnJ0a19pcHuqJnRJfnXiyGmLcXJ5eCBOfSZIEM0uBwB8r/Qnbzy
n9I1k9kIC2nb5Zb6gB8UKIix60MnwACdn4jG8L9k2ko7evySy0sQVM6eHqHlu5/NrQFWef0BPmiH
pdSGyHugK5NuwEiJmV4Qhejc8ryt+nC5ug7D1BM2vZ66IFy7IgLHo0lnLrOpQSlDNydn15z3Guog
RU5Rb2LHgCzzDOPsi8JrFRfJoPHR1vD6Uz8BdlgDyssCq/7FdXQmCSBiku/MD1FZIRjcXUp3vqCj
ccba1PtDVGH0Ry1IdDKhSXeOKxgrzPhEkeWalJpM+Qxemm7wZhLxH8Ax0/Li7xq5bM5FZNkalpOg
kmNAeY4YE/98j6yaf5hItBz//UUjFtGPzhXSbsl7UAEQAe9i6oNfMqc+xnojH9q0mC8OH23IAa9v
KjLPkpgyLdJ1uqjUdUKMJ2TSdlXauSnv2bJ5E/xjvomvKS2LoUmm/JUWISAVPAxIHeYvL3k2ilXB
d0chWwBSBaCSqhqayxIq9HcIk2YG7fcc0NcXX7bxACoOw5Aa+58NWkwrbF74uXSWkKmmnQo98TTD
AUtYXsN9PYKjO2V4PF8VHAuHjCb8cLxFWVuMrw0tn7hq1Gd53hO5pLN5BD8B5tsGLYKEOcq+MvGW
/LIpB2Z0DG+eJPatylHtZJX4R/xSD6wl5AX1fPrEDULJz1yTVUTeN5Sl7XWyfSNh7RwiYlcMHixs
LUONWBKxwJ0MBZiio/LFlnc1zLM8Fo9chIhiZfrh5kLcpuNEGN+9NODgSitU9IWW6k+Fwl12ic9H
EC6BKT4tzNcos13tWmNIiVS0tGH4xCtvpflzRislSTKqIDP3S4WOC0NROvCwatPWCFUTCaWqPMOQ
64iz7ngZ6FJjumUHVhua3gMxi6My5/0FYdHW5NqppzI0DHaOBWBebXhQr0knnffIB7YgaArGhKpl
whWWefKYEcTcvcJcwbI8JDWCBmetl8EyFnNo69Yqr2qp2hjJ7zl4sC/wh0qinlVvvtEKsc+Nyg4q
AN9IP8b4u8Vfoxcjbm9+J+eTBzpTmlG+GI41g44SKbpYr/hwItP8jw4Ao6HfVw9h9qFEDP0+f++C
AjEFi3ZAreaScFQIGXGdGyT6CNYIzJ/7xqZ+e7Rhuk3W0JdiRDvrqg8nlFy3bGnXIL865U2QvZND
WepsNMmjo1yGZsA0T8lY1efjZ0PY36dLLkZqbBkEQe0V6rZrXe/gozz7brxmsXt4kujFkI1cGJXh
bAa9merhW/uocprWJq/NpdYt7SEY5iOM/JHK+uN1euRiVLbs7jGhG41tDor5EoLTpY503awNNDPT
NnvZKaKisPAxv05SYtQ9rybj1Ifsmi2Kb7aYxnFOVBkam/m3H/jGocMvdJkO+2HBM4KyIe0C6p4x
GVyPZX4JiRuZm1p6wm/lRA+PWI7NQ/b7/E6FW1eY4/O/NsdMTmN5BGf5muq0ABZN4JfFOaN4cXFZ
q6Ziim2QD32ScAkE5isUnja12FbavAx63UOJi1VXRx3AGZMNcSkXAeyortI9YlKpz3uhBj2z5DYl
1hsN0Be9ss7qkXhU4gTJV8M2r9rvvP/5inGi2Ix93gCSW6kPyYhgsINf7bAEMD0jdDnpNYLY+QvY
7Xxhkiv47EMGXKlZ7AgTVWYX2o4AaabSwZXiE7l8ewcfbsgvtyIMGOk3jsBHuZkSAHQbZhklbazx
dCOAQ0LwzX66UhSTfdMnfOXz58vi3E3UC0bqeIdfx7xG1gzig4SjYws/CnCiP1v+4FKwXE2LZ7IA
N7kP10koHDybvoVAlQCIHL7kHfVitxGdynPKr8Sp8QcLLjmzmlNyjVg6LuUgfST4nJusHUdQk+S5
O+T47+1guiKS1rAv7eXVj/CXKTSxMc5GnllTaYE9K5JnzIIlQkiNO1LZQ6W/zRCpnEchq5DQ85n2
ygYIbN/vVS/+S4slAt5Tu7+7sqyeSgGFitjQ0sOOA3cgsEFBGu9HzIzfl+/C2JTtv2jEmz0JauG/
9DtVFk1VuS4iNmVAMKArIFtDsD10Fmz9f6CluCfFQugnVNs/ehjYQpVsFjFwFR+c/M4koZKCt22F
ugksN1kIWCcyZQNjyDBn4mvtFFyZa2XbkZveMHdOQcJSGqHNfHS8vIQtktts5eUmcfvbAU2GF3JN
cSvrzw6HHWwS85By6Esx62IOBPD5hju/FmP28AnocJo4erKvTE7qh+Nfij/XyyStclrc/gmO8wC5
V416cnG9Bud2qIc7r07izVyM8J5/xSVBPN6rfLZu/RHMNoHYqoGAC3WR4vUoAEilYhAnLBsH1xso
1dSl9FuighmFPJK4FsbldjN1pNfYZr9UrvXXPsRaDyeuKh/NURPrgWzUhdy7hjfLIwepADFBIWCy
wSm1TKo4cRWv6bW0zxriyoVzfuI4i1Q3XvmT4KMkW0ipndRjx6jU0h5o2giZHd0NyxAeRdxpNZ8i
xHMPsCaL8N6G0ZNP2VFW2bwvjgRmlHEdoLPCgnM88t81ZMdHScpp03agJexKsheB27FMuM2K/ick
zbcqspIQw7Cw6btd+uaK34BImwMkr6rqZJn1n5z7DvOzu2txiip2i6SzF0luYvB8MQPr2giqimDo
CUKyZBZsCQwTc64y31mLiSplGFQrvemIGowtaVwUDSATlK+PK6F+ZQPXCnk6LbMVhA8XrxsKzZiW
hb2GWzsRGw110COFLgcEYrkV3k3M0exVaJyDwSZSfZmAP/UxcuBE5SwrOzEm4WWzJeZhnPqtuvsJ
Ksx+ImkFePvszA5/YVYGMeWyxBHFNRU45wngvhWA5gwKEcQ5m5C8mCAuagxXTfre/oZkKDJUAWHX
iypRXxDjioxotQiKKIWHm0QYKZYo8N8mE948zADByaHGA7WhJOMre23I/MBg49J3SO4qQ+rb34zl
1u7c05c2QzfuqWs2Jht4N8z/jOtTxxb5sOzo3ylNvH0ns++ckOc2EqmEogYA/m4juwVewh3gm2Ya
XfoELw7EgNGF1diE/qzy3bqK3bwY71B1/SGKL7GDPo05N0hg/57kniBkbKcsG0Jnb/G6W6K8WtXZ
+yTtnCcVEZq0TP5zfwBD29a/9txSR8xQ9nrW8x/p1GwMIbeleHL3kkP56N3qwPsWZfdiGh6dzUGq
SjnhJoLxNChDZ6dcg7f8lvF2zMwJURD3ZJLl7PpiFTKX275SSYXjzPxeAImFHna0Afs+aT62jk5P
HHOsMCLWh4NjezHdS05ET0SsLxdERyjjld7qExM3ZIK62a5KDwQgg9aG8eqqa+JD5bATlrH41ViR
sqasqdfBToRrlwp6jp7dahaivDRn1y65+BwP+028c/ff+deqM7B2F8TeIjqAIXeaUub2hmV5VBDI
RN22VAC8SMELlnTZsw3yurCm/5q2SGSZHMVeaVX+42kVU/HhZVy0NLxxb2G2Kor3Mwf6f+xMK6c2
fWRnVYr5wRevluvVkIWOTCmYsviZ8+7+1rO93Pjoz92O+NQgOXxwdndAU3/ufwWKa2sS+AkVrkp/
U1Nxhsoy2IAtrtOr6yUxFndzITWgXpF2JTn5wglvkMzW4WFkWJHCFlc/MYGf/f3cNoQVu+++tnDO
bl7sEtBuAQ2xovyawbvFdlkWlMhQiBNS8dcveVLg9Bu+QLyvtUTLz2vmUZEANORQ7mrhLoP7fvRe
zO6eQQANNHxQXZcguE4a//z0ua7fGH+/Pr1L69EjdlmgwGUyVHKTRPJQpQzj21sk2BRYwjpo7TOR
SSjFniTJF4WdmTx9MpUrVr1ruFnXxFdbhRzjGOSi8Wp4eRqwlN+rvItUrR38oDy65Ogfaj7T+6Bb
+eWKd/xrvt1P+oJxxwaxcI5bukk/4h4G7kM7Zzrab62yovFCQ4k5TIlJNx9/fF2z+NzYaKsk3V0M
Kr+lnFFlGA27zKnVxKdDSZgAG6meyC02MpKum+4+e9TcKQV93hLotI5amMW0LQsQyaGPwYN69rDy
pR5D3RMyiW7VWRkcbUMXkXLf9KNYI0P4nXvX/2taEbAz1l+9UWDOfYG0aY4WvaTTs2wQ/+6ZBrSI
BKyBXqF8I8yglKMY/VXGIACI3QG+0bzfgBbLQHNI5EitUHAfJVYiPg81stullKh4pBaIovYXGNmQ
LHuZHbQeyD0guEWG//59BeMSCdpPW8Me/+moJblNM/JDFelB69dkZ0gUf4E0X5f74+7s7UC+g2FB
e3gttn2ckJ/GPjCNk/GI2Fn+6vfPHZAKQo8r9tuN+2WeblVx5s2d2NaKMUWvDKk0NUzW8eXwq0rz
s0zjO0fRiRCp917ifvfJ6tadbgJ92VKjkJ2+KJMLkN6nD9iCPIMx+YDI3vp6+ClWAY3NEtl12kPr
5BbH47pHxNw7aXnvw8oAgQwmjXOzI2StxrfMsHPr71EffgAKWL9JnuybbKeXGnTC0SWAGjWr848b
e6cMszldHt5ijY00bF1tBf5kkV9EgPRySn0fvqtzDxeS1XOSIdTk4KbnBHZ7vD+4vr+yGxHXS+Nk
hjc36AG2/O4t+KQK8nCpM+G8064uNLNzH/0EKfZgbYk94p4zjIuE9f0fHWBNIXSQ/5Q2t0z8wbvn
d3GmGqYjkrTgnEWcpLp1AjhS1syiy4n3NE+HSrh+vb50A9bNCyQnLmB/5Xbl+lCRsHX0dRmRuE8e
VWZLcB1kYApuRcbdneJClYr8GThQTvFTWlTYK0oCnuVPGS+0wgCr6NxILKBZDarumk+oobDbyNcs
9PsIL2papmd+f80km3dChvYXMs1R9Lorn0EBKSjWKbsy/ze7C2mtvo1+9W9DH+V4RgdtHSLTj4w5
Fg3sAAUMQ5QHLtbvO8+Ah3oV461gd1CE5urahf4K+C+wlk1uyAG+j+at3qaV6BRRA1npXEk6f4eb
2rK2/gV34r4AQ4DXPxIGr2q698Hzs/p1wZjxgcdlUkm+4ifhGhYAySt0GOfGGSquyXABWLwwFE/I
wvQELPa6XFE/ydZBIehzZshZXKqzxMSFbV2teM5dzdbY+ofE0PVV3d5jVeTMcN7NRsbrJStp2j53
PDDPr/pghi4wS3WMkdUTxYuuBQ1QqxMDNWDsTDG+6V9n8WqSEf5Ln/9pVG2RBscQKREVhNlzJthT
GaWYuiTP8xEFPtxavlIL3GMdSN/2ARjvlf+SwMtu2YsXPAopGt5ROdJfRNIBs0tTJU8ugtq29nPQ
mNhlk2FV40H1TFcKo09NOFC4xwaVoP+vSmugrwuuRJGoCr8ZivYr2d9XCS/zQGocLWMyFQYlGIov
Y9Vxd4McIVssTYf7BI77FN6eAgJAYDYz0epqpHby3SxpmdM5l2ala4C6kcA1fRtFU+o47EmTJBbL
xGJV10ayWQdrBTr9n8ttuFLgxJnz8t4djVSkp+sFA+h1a9qehPJfs9s7ZIT/yROdbIfMUAxOykrq
9JuK4mvlNcY6XLJFZ28eV7WYdblD48+2rsPOOd8/c+t6UfzA9IzJXNon0s8BPbIYygdjk3/90nWS
BKKf0jAnJkWptvPiAIhuH/1xwYddZ6Qa9M+uqLc86IeSmzy91NmnVtugUHtgXidc46syzIxMXsM7
HW6QgTZNgSHh5IQTqWlnNtXziA3iDD67/dheqvYnR4m2oUQK1t6D4FcV/LCaEOm/YDlDXrFQJf+J
GRL938zwwuQassjOhAuwC/EfmuqqXo3BSgcdhOJXgSiDzGCpxgFdExuEwBcXmD2bbzo98V3CVSeM
BnzhmTqD4xoU6UNLio0wlubuj2a1J1bIleuAkfFnuXAoc9PRTWa7ARCUUr4Afyl1NqSr1DF/SxlF
iDC0bOjkRcuDdT1AVKumg9R7q8F03fgvkurCTD4EpyX91SZZuyF52rp+twOvnmf407MWRgx57al8
+4MSRWf4bG14Tw2138ZWw5W6pPJHVKtDoJ044CVdm13AItqWr7bObn+ROCGFdEugHpeshiYp5hXD
F+8ZI9AKCEbiqpPfAC74tdq1JCv25ZQ4qpv8nVBmTorrazxfKWg38dgAT6ROpDFAomyKJA6VhS2L
rEpLCoeOxrVbyWS1VUc4iwIeIJrNVPNCpJKJLH8BceGkempkRAoR6AZkIDijKvwGNJwJMPE8+bPk
VXUz1JtGY2aKZmp5VF/kmhWXpyHwg8JRMsi9z+j1mkLU9EHooJi1h84G9xfSa4XRPK9dIkYqMCvd
ewVyZ+t9ZuKn7HTQZK+QUpqjhMCDdNvA+wmor2rrXw/095fg6OBugeGTGDJkqhv0T/kHBNT8pUKp
qeShNeOjOZvv7KooR/vQ5VNuzT/8uZp2/SQxh2AnF5r4jg/0HWExX6rjfI8cab+bFLEgNWvDPbBp
PExx/LIf3XuH4NwJ76+EG73bFqk40irALfov7cdrDQxGlaiDxt6d9nv8l+r3OYGnuBzPm3jmEJys
proj4DKoKjvBSIPZhw1aRDqEGi+UzBog3jABYsSOn+jI28932hpxWZaNb6bZDGnYXHRNkG7bqjGm
5Q62qvE+IQxMeE1/FRHfCpYzhV2EbqAr0X2c275TvsemmwrISgaIWC3dFxAgXi5jUWXlqUFDKwN4
QJFiNJar8R/VA6ye+DIP9CNDyVaXi398A25x0M1wT7TQnXI4AppO0xluEB0dm/u6H7+0NslBxMpB
quV0jMkxEE9cPLS4XHQb1tLayy4Xt+YzYkOekpl3ya+HTR4sPtf3DKBnhw2UJtTexwFhOyQm1OoI
lJChCnWci4T8KiApUl+ummrMOVWQY8C8FfS1dXBU28U+PP0BbfdDjdR5ijAb/5Usr+xbG5ZWRL6l
re+cKw1fop+Zwh0tYmFCDkm+6YoWsaHwKAKNpj7r9zEdD6KETnV6U/xCSFzEtOQE6SyM/himi6/7
chYt0i1swTXQM1erGOSsoppl0cZ34NWUDAOGoWAMYoxXHAVC9XhEubbdHgKniC8PySgtH1iSZTAc
Op8oEwox0M8ShRMKB/0OrLcyFs4tJagnjzxYH6LWB2zQVDW/dlFFhzsQexhtO5CqReNoaQPvG77K
KAQB0q666TMjrXuG/dGJY/LBuxzYiFrtYtaPcFS8XMohN7AaYU82bAGACI2QJ501i6GYwLUZhsWR
AomuUkBNqZGQUDLbfVmF3TYSwPkgMKYRSSE0EEi5sPGMmgwAsUc/GwePqT1/g7eZjyYgcbsj3Kq9
etq71iyBAk5GQOjJ9zmQZtm56Sq96EMCeacwRuEkKqM5Lqe1vb2RWF3Ibe0tM6G4jxXVpYaLst6K
k2xx26mBB15VDkELnegz5nPxVPBtbaSRsIrNqsbbSe0FjCR9nTml+YUw9flMgWh8h5YxwQxrCdvF
Dhm+HRewoQAXuLiUwjI6WjOad4rL1kCpNRjYbr1I2D9QxF9uLE0KW97HYZDdoFQCsU+XZ4jKhMn/
KAIj2YQNXLX0ZRdGgPwX1n0JfXeNJNt/P2WJ75o6t62Hx7Zu6WsDO+rE0R9akZVi7drAz6hq5fz+
pVsYCTN4qqaoYYlBi0ZqRQBMHr8jtqHqjRPBbjIfHcpUWUX5sE9HHneJ8P5w1MQdx90ZeCHmgaXA
0dh72jnxiYOwDCOIgaITr1mlJx2Ihgo+TS50MxXocmFnW0xWSnNkXdDbEO1uvAqWyoziT8rBviZQ
Vkh+76TYbc5Eep//mIL22sxGRr5K0yUeFLPllWPFwhDm3wo3W6Xr0eRKC//Ovq58ZwgBmuFm/jxE
6JHsiNkXrQ+ew214RlnV5WZAMktdC+YKtvWNvL+Rm4VK/XsYfICEGdRq59NE/NpJtT5ickU3/hph
gtwxHs7WsmS048pswiOGix9aShf2Rgg+hSW/zUxX/11pYD7+N0SFreT5tSxcXUV+TDArtfnhtHAy
mdgTAJZ6JNvv0LtRWXfnMNbOuxVpW1/rVWmiAE+wXHi0eDMeOrL6AKnCmaTugQ3dR63BD6uuZoBW
vaJF6WjCsrBTcdW7LqRkg11yjeJ6SmQtHA4vmWanWKIP0XreDe4WPzaI9vPkULuGGR1YVCVhBAkv
pujgTb/RB+mPTA7iV86Df3LNVhUivQn58uANAFcshkG48KSheQRXesQvJB9jnPO8CUrxJvW+PjWz
38Y194B4rpGroFyBadtFfuTuydo5lSRN0Jkooq7Gss7gWOPNAjEdCpqfdGXb8mkclV/jkhwi2wVt
d5XOYbXMy2MJ90qe4M/WU/4i/Fk4I8t7M/XXwqocWMVTO+xfybIkwJRGNl5wPXkWmYxnN+5ddZu1
Dlf55R1ukZAMuVnHUBRMkO4bC8sLqiRuapXWimMBxVUioPaVL+BKwC0dhKnHBvbTmiN3e0cU8IaJ
bb8PaKfTxJZDh3B+50HKrJy/i6OY+HbRMvbOAgmPtPhro09kCFQ62Jiw8dSdANaR2JOPGpSFLbFa
+c7H1eyhiyUqmZ1uhlxXzMAoWgYJEccS6qiHdRxQWWtGct3vQghBcHHTUYhgMh5zk6zfL7eVJk9Q
98U6HDH3aCAy+uf1WOTnKJMWAdAmry4lTdQ5s3Lw+fXApnlFzL2I2orShlLNBA1huYKMa0BP3jnB
JhyyFi29+8Ag7USOniSoDAC9g1IMzQ2QCjt6cJuHGV7/MBjae7utICK0dzM0RVxz0EE53zD4R+Uc
tcyhv18ZxvIAe9LcqwTUUu0LAGYrGdOMkaxVj5Eqs38nwhs2q614rGhTm48IoOJEbmac1vK/Xtb4
jC97K3Vqfk0Y4OdxdHeXExc4IHLyKoqn8R0Jujn+nIzzZjbJOp8y2x2q9scIrWHAdM5wZ1bPQsb+
RDRv1AIWIIbF2gPC/FrUPkp/QhqA6uQgs2mUTFlN2KopKPcP0WZgVHPmH/g0kKtVfqeyfSNYPuow
rtGbU15alJ3snILGcNxYYqcVeBzFwlcUj6KaqZj2TZj9QbNMF72kQR9+LA8zZc9S3jEW2Xi3eXDw
BuUmbwGlx5HMaGFOwi+CJ38+VE6wVQgMtGKzrYYcB70uA8i70/qtkrANb+LoImmkYUCRzrUKhP1b
82Mmmd45F2c9x0nF8GI5Ue8/MuDnZIDD9v8lZvDt8AEJAfnM7SE9cO7/Hvx24c37SXTJ8jvC16IZ
fKD38KFtzJ5vV9KyB2MlDes9bauVtPmEqhweLhUsifRtsTkYcn9BrSfB/G/3eUiWmQFIINdgb+Q8
9hDoGMeppg1A+ZVWNaqc3Jlu60P/F744xoReGAoW1ZjiJA8jziKMzLzrOzHPe8Fc0xwoZxJSPffx
haIfN+VIXnE4OClHSOztL6Us1Y6Dtr0P5CBypTBdRYFhNXGRLBf5TDD2qUxVyCfSeqlexLHhMxlE
j273tE6sI3LZFcramKYTlud4NlFF6S1SwGOxmBVrBxGgV2VK6HGY/sh4lO3v4rWV3gmTnjSbFjlh
jqBLz5HaUM42DJLMb+jq3DdEW3z3k8ZZ0iUMS679ONZePdmkHOzAhrJwITNw/jKkJWWaqlVd0Ewy
kzNsdbCJ4AOAxhHHPZ+HhPyppxdg8be9goRtyjy8P++qRzNVuEfAOMwPpZxWkTy5HfXgG3XLiLbF
M+KQlWPYhKcLiWji/x9gxUtCI9JzqJtyUijsMpGCPdWlD2oFxcsi0M2nDJ+RPQnCCobfCM79JkWw
wHQImGFrdHvBP3gJfhj8flq/O5fCpqH6Av/lXKpUfxB+9gvKeZDoO66w8mLBzBcGtf4OFWLbghoY
0XiAQ1zIyZ0mNN+cCOYDnUW24zjg+F/TRVMtAkgmSs3OahV1elduMmm6ofQ2iZokhR9iJ2u/8Zjw
LePbQWe91YNNzl+84589N1N86Q8SRwUKU3H/3q5XVQ3/9ZqxMu5OnLc3tcteRogy8wcuwfMJUL7q
UktL0ScgnFZTkBAEQtrcn6P7jGNNx5G1XeGJ6lt1oAWRg6JhCP8zJGk50Eg8DoN7XyYZ9KdvsuM5
xxEo/Z7xyRRhcgfZS4kJpTpqg8tMBLSgPHXst9BA/AmPXiRFpWFiX+41WECuJ0hYDVoKXC8+t/+x
/KdPnANaCqm6OqRinba2/fyaMjxj6tNazTklkcctH9tkUzKQqYST+VY1vw5twDd/9vA0HDsLmDUX
afMgn+svS4vu2KAYBBi/fdjj/27vdiHmVV1MWy7hthnoVnwbSMKtVXIKiTpwx9C9aSPbeTWCya50
8UNc7riwOtw8GXZkbGnx1QiU2TNwE+n9uHTH2z3j50TroFnMp+w9agPI9rVHGOI2A2woXL09YWn/
EIspdnBHFMLXPquloKCkAok1Z2w4B8vn/oJ27wDhaabUnJEVbHn9Wao7lDkj6yVL8CFA9QYOi6U7
foBjRCNHvBPOpIBv1IAN0uCVFEEXAfcroXDH4s5ZoDW2lxF185UW2hVPlAoJKGBmpUObToWsQt/1
zZIquIbTqrLCTlPlEAhwuJ6+eVKIco7PWToxU0iTOr1Hk7QDLuDys8EIguwxqtZNmeXews3Y28os
eH9Jl97il5v8sMlll4qNjuMXOArV7cFcDicgZ/TvsL5usVIuvzCRFuSEsYSOZbLZXJCqTUWrORLW
hm47ADWvvGeCjr26nWptsLmin0ElpxD/2S0s5/tVhv3AGakFovBJqEUgmZXAoUaNrTINAd+4ZO8L
oswUviyv/AKGKwbjYc5WQOswKqxOAHzYirFD/5UQoCUccxAk+Fi+TqmQyZYcZOMFAIgyav7uPs6l
LRefEBvhrjGAQqzQtBfmAh3du6Hbu1ZE4iSJyKbP+S6ndmQBuCSM0i1/o7DUx3WSzclcBOF7dOI6
xGGVPDVIDjbWlTx3xNwOxtehW3Vnt6cOfKiHcuTrOFJuJLNgIF4Wf0Fr/Zr33QYxymiDGYMhXfDs
+ZeEURHUZ6QOgjxfIn3PTwXQW/YPlNw/eErzUzu+pJkqyVBp5qJ/TKmJuZzrbsdclywripwtCQI7
W2WmpJF2yERTVg/4JqBfJ9C7QnDhWRPAo4vX7mYPgCnPu+C8pQ5AU+Him+MyTRSskIaJWu4hH0MT
ZGIts4CY1zI2PMEub5CQOB+FiyAOTgnRV2c+c7vfdvHJb0U7CvYaMnKpmp+YAB+R22CdhPTVT75q
W5RUgSPuayNAowCajXeR1Y3VIQgfhx0kI0BgtUmN9U2b1z0zc+HADXD6Re6l3JIKXYsH2tSThfLC
z3HJL1jZs4/Eh3ARl+UrGbFRyJmQpQUhByk08DVElNJ3VMA3Zp7L3hDhFo9GbMQiUEI5qBTEqbCa
O2ELqwDevTCKFHF25qeSrQ+s4toEHdy19KhFql+bOSRE6EyM5NsdYU7Q9AsDLYGTm7ZCR2kcHbvU
11J5taF3CSmEwpdAPCvE5xuC4mIW/DLSh1LEG3ZcTeEUZQrr88fYh7V+Mr78oVf6n2m72E4FvITz
mN3EjK7wPC66EbQ4lKxNsRuakCxf1R65PNTyAOs9SAIv2dmjF9mJ0odgzGt2LKPWYqi48MiXyjOE
7sRI+Lb8mq15fUFOfl7us7j+5SnWQ54r8y8Hl1DVglqMLHGiRZdyAuZLwp82GFKciNK2MRcwyAH0
zE33nxL0e6KyHyuIyFOLhNQhHnpbO4SIsRqR9F1SF4JvXbtfzY5aRIByCJ/6awQCmbumhHqLMEKM
l2o7YIWddb/nbxlu1YSY+B1HzWi3TQ/RrdGgAF/TpopzzX+5kV2gU//4bsKYoANxdmJZZHSOOJHW
GUmOd580uXw/go5gpIER5JLmvFpAmk5x5GOCNhfftwmdc/jbIrO8MZVZUluCAQo0fJDh2ETDGZjv
sM+iHazGbDEnPGLE0ERvmIZ+/z4gZPJzPGOk0VhX5r4EDOdm8j2zSTJ848YSgZXj6yXJ6z6EWfZx
qocQkKCooFrieoAxPZca+U15gipNnnIf8GUFSiKuXIuqwvfd243RYMTbRyq2mNNlB9T9YpiKVQhb
N17y2dct4FblHbCmPcyb1wvhRpMeuWg51YnKUSxixN0G0pZ4ckYxstCNy9VBnsailFRRiK4R5jNO
RM+YsAR75g7kKIguPwB6T0lZ5j670Su+JiGpTFS0UZKafW8Yvys/TJVxyH6mN1TNxkgaQx+ZxqPH
GnVKqdxLjHTzF97Eqwkm5qT63V0pLRzfEu125lVrGeY+Xe7RqurlyqaPt8A2GFaSEkPfRnC0yzbX
6tP5xrV7g5k2ahEs2wYQGjzXd65waUk6hslIt8CK6lNOkE0OA1U5cbaupFrx0uhAz7Sh4QQEVSI9
PSrDhAqOSjnhcmMRg0PgoHpgVxk8MyDZEuQIYDzkorQ3uBEa5OUS3IzSvVEvlcOuxGoFz8NuJps+
DXDyIYwwWM8CEHxySncfb5RX+qAkoWLbrkk3pQbwQZfNdAJ5klrwKCoGMEu/h3Anc20uGsP/tkBY
6vyA2T4SQ5C4MwyN7sHpiuqj87PvQgposx4LJiEfdV9U1BRbTd1Ewmf/UGarN3lZa62eVUBblzTQ
THHAaEsYHbOae4+EsHhtxV7gnYqK8WJuYdWgJrVwy7SQ+6Cfz1zHpWOj36Ir8xJp65qsHKsANiuO
20OvtCPYEG0mI+F2r+lPI5CpK2eqiCm5dEwjR2hYMJqHjcN6w0MinEheX5yhVEcGlKMxvJNicGV6
0aPM5KvGLF/xnNiNhZHQJC2kDRDdb3H9KKbNKOiGjoTJJ5l7hV1ux/y4++gt080Y/9Tti5oI3bK+
iMtk95CqXkpcvn15jV9tfOHFkE3qkSFEd4ZRqYrk6pDcJ70SLO5sGYqbEb1uzl7pRS+oNr569fmf
eE7UPLSqUjbIDY7HbkDuCcgiRKgT5OVqoOYueGFfNmDDkUjRwOUjfbH5J/Ct5DelO2QU2emO+MwX
aypkXCXjuG+WgGSxnWlkhQjnD4iZ6RItVCVCWmhpR3xqsELgP+vB2fWp+knP8WgDOfBZACw0RG17
47Rz+MFsYwG9MXChLlfFAXHre7pkH/x/ASLFmmOEmtBhKWoCnJ6NFQT/BflKrCA7M10/cqeRYqGS
3zD3aYdaVjTjCRKEll4mr1807rMPvEr2KGsAYtKjG7VWPzuKcW5s2OQ30yPfr590sff+F+6/hOZt
bdsqtexsa5u8D99rkM0r99ypeN7u9KwFqJq0QlabEHycngijKmyXQPJPLM6NVKBliPGX+XG1aQIW
VTV1B136uNWx+KUMIYI4tidPFjtoO+2Hm/GYryXr2Xgzjnc7KUrSfzrKZBsB4O0tShG8ABPWx6Xx
EJ0lA2zC5fNMrRde9BVCviha5gA5TWj90F1RXe015pc8xgMc9thsJKzbJ7UIwzP/Z6gkbLfduIo0
WA+NH7WzDYNONYIkcLisbZj+GARL/oAGd9bMASiRxid/OXi6SIry9DzhDZgqoKQWlrFcjO0KzjLB
8/uIY+FZKKGxcEILhRey/KdT1HOhEv1LXVWQZ17qwmq8C/NER8EucZKPrhMZH4jYFNqAZyqeht7M
MKDyL33FhXJJlB/B8ViDjdB1ELmYyl5mOwZyeXH0ymMJqRs3Xk+I5Pc/hlXdjlL1x7pxJmYUOs3q
4o+Ca/RO+VeZ3fCIjcIFS60MihgXoJBv2aoe0vnHMDtDAryLnd0RHSR9omMS+geMh2U06xNZHwFK
DioLX1D5EoJ6TbhzvJiLWB4UvmZzPf6+3nPTIMi2E8z9aQOqF3p0PV/9nFmOu2oEnYG5l3ELxpY/
AtG16/BTjh8RH1yvLvkYawDFkapHiGh9cpWwGB6SHabtqR8wrEUKYjLeE1i74LfhtJUHqgrUP5VC
wqTtR1Abxz14CWsBan1mPtgRBvHIgl5PapjQ3tjLteKNeUeQ3m6SmUzNSapoTtvoHKHzJfQLdtdG
PNnAYn50QH933bMXSW5o/SjLMazrvdL+aviwehQCHYy3P1M2BSsgjmfEGXF6pSJB6lE6bPbaKChD
KUtyPcodXHKyztscbTYHG3HGvGu24NP0T2NDsQOmSJBhxul9jYo5gEZu5MsWWNsWtCdn5mZPKX1B
ZNSMg4AfpcPItO6wWhAU6ia+FppqbSDFsvFhvkDnFo2Zdow0ojT0CRh5imSsNMPzF8spNUsJxH9g
axdBZQAr6BK7TLFF5CF4wzP0FdfCRIS5y6eZr67JLmIC3ZoF8VL6/aM5tX0d5B2f2prBrIBp9lbA
3NVIdTbPmiLwc7uct2lRygnBwmTGtpitqWJFx0JwlwjA/9dUZ3YoBxXPBTso1yhKjp6az1AQaz6M
PsNgKg/SslLlDIkURGzt5FjSdnG9Ycb5cw1vGGCcFx//Q8x39VEgG+N/eeTL5GgsuEAltXBYJinb
WsgRGtJgy1yY4xfX/r4Adru2EjBu8jBTq1OOGFak4tbgCs49Oh23IW1+LM+JdZ9f1kp9kuN1o3aN
moUJaFmsZ8QK1fHyH7qH2/9OL34dOXV19C6TuVQMGTSlK4IBFNby3SxPLPLZXaAuhyBBfvNv4RjZ
/uQBTQ9YuzTx/LUzzuz9CgGApukODRmhJ0lJ1IIiMYHhtHN6luWdGLZlZKAbea1zeiersYJjDpZ9
41pg7o+yK0uBFi/hxxACne6r8iKExcF95k1aMHnNZdsSFMgZJ7XC0nBSH2P8BDA9Gm0/E3eH/81q
mubA90vcAazYITR1E2GAJMwuL4HejuqLpTgXoLQDrXhyBS/jZyHE71qqOLNCw1Eg0B962NgQ1Lwz
bvnydGYphAEOcfyt0tYN1APn4jfxIB0Sr48XrHXtJ8bmZjZUXMRBZ2qcNXe/eFMkSAxrqbM98k+k
htUULdshIDdlN+TTEKwTxumqiQWN+cTV8XIJq9USmJ8RaUkpvMGbVwQFKRAlEHceTlCYLeTmhcx5
RI+SQsHp2VeRKF6nqtICsOOzf0YNb530FHvT9jdCfbjR9wegvlZaECW9nJd2s1mjoAtHJtMwK/TK
cXq/Rob6iDzKW9gfD7H68DX21trq8gJb/e9d6eYu9Uhq7wbK0TWDee6WRRSAXV2NK0xhhb4C6l+k
h97vQlGaNhO9MS3KktczLmxfv26Ksqhf8x5JzqjiBGhnwSLprmMp63No6jBr6yOumKiOendKsvdM
pu4fIBth9K4pLNnOZ2NInoVqZGdvdflh+lTVW4acPQ4zp3N/CdxFKXIsvwa+0Rvmi8kjUvymUynu
bjMmeP6OIkKRNeiJZGHzLtyNTq75dI0QLT0Wn8OcIBSxhVVhI4VRHM6eRDztf9LJ1+2eelGKGtN6
8BoRtLVYDBVG0J62JULJwZTb2/PNmHGOa5RyRKDZXv/GCNPyGzXHHZaZFuMab9/uDGCEuL6xgHmd
ZWhv2z8okth7nl07vFAWEyLClMBSGBzH0BiJmYGbidlKzxF0xrZfOU7ApFdEeaDbhkm6mNzrcN22
LW+fVHKpOTkPSJ40lKgNj+vKYDKKpFTa2yCfRK/HDfRL79/YzO1SwJNS80rIDe/eCyiSosNEmKdW
Bq8p0vdrpVttY6Lx7+N/GKCAS9uVFQsPPPMHfo3o7vKIVi4OHMX+nQhJuDeDAxpvbEKqwN9pW5qk
DH6z4F80YQ3OwjYb6Wg1oHx9TqrTi6bFr9cJerzxP1WljKCc6H15HxvFLOZ5+QTe0xUGnKlBJHYz
/z5XsvWO7j9+pmwd1SSbxLddmbFO6rXoVgaOqyi+mrVJOz6UAqHi163dJ2fZb/daoUMVHQXvgBVu
x5KH7f4Ntp8inbr/q4ZlmkG0V+XZ7mOMcr7gbp0QqylCT1MF1Sjke7aAjkxV4gJycGo5WTAv7F2Q
LwxYp3XEmFTQJcAypyeSJ1mOW/Ityd8RnfudYsRo7FKQ15dKhwkIDpUHT43lqm8Oywjkvf90yCDF
yyF3Vz12QQgtg9aKzEz86/OAWg1CBLcqyO+qmdyKQsZOJzPvoRMWADgjQIfgxomtEdAKWVv2ACvO
96iDotyOxtFlo/8P0wym1UKYdvDYrpXtr1GrKwr0MnK44k+PlZDu+HD+Iwq95rDHj+O9JF/EblNP
KcK9CzG98vLKHf0GYFHtmEYM95n9R3/zLj6eEF+Fjv91vaQuPAXctA9Y2fiKlW+5B++nnRzAe3DG
RdSB9X9sJSB9sTg3UfMPdBpIM2SbFRYmAnivXB2bUpzP97juWW67RoSiOdCVIyyCGZ+sBrLPXt/X
Z1aOwTKfaTtJH/Y89c8V6fLhVnblUt7u+H7keQCDInvdwgj0rHh8NTPi3PMPruIwN1h1yXk2Si/h
tWxqPPphrzpiRqQVSC+rRPnaRr4LUhxJfIv33OmfLF/K6L5hXUKdqOOTrB1xqbfnw7lyJchabdEk
Em7iQ6s0S29l+h+dNM80rNd5zsl1f4ZmdX6GaOrqkp/9JSsB/w3QrlGyOPFIKGH4NjIzDZB8oNMC
hB3n0ZAHcOvyJSDU0ictNj+DkNuRF5rlhW7MQhuf+a+gwcaZ43ESNUaO4RBKUQIm3fiKLUTiEwnu
H6Md/YgPJM4HxI00CwPr7vJPQIDg6fFLak0vJ481EB0IXz53JY1qYoFVrSroB6DUHoQn6IELMGdw
KUsOx6tHwVhbebh8F5ipmlmT/4gSXtFpSkMle7UDi62un6i3/ePCYeHXhF4NrBFQxNTXWIfAT8/g
d+O+Tbj2vzc1D+EyJRAim1WmX8DnofdBcrKo/eQjXatAdzFwCE5+s94QhNEWjtBBm+3dCkyL2x11
Y5E56hJN2keMEeN0j00UZyK9g3Yd55iKxVoxZnI5xgz2QIgymzya8mSweG1zS94+6/DIW0W+VnFN
4eIkhesQFhocSP7DM85h2+ivglhaZdgBeyjpw8OgV0GKSJDpAbT6Q0E6fu/FS5/Hp/RNevK2S0r0
Gcq9C13SjFUsUXJrcmGKNBtv0eDJJW51iQcJ3Atxvkdnceuc3h+gUucDLXJ+LeAJsyrByEA3fAuL
VgnkJ2yhHRYQ7PBKbpL6JNnc6HuqYpFgb53VRh/jQ/nn2PfglHvbjCO+uR4hz9n193kk/1gSfUYg
14NlSAdmsZsvWQVaaVkLPcoU4O6YL5dK7enhz0+Ihyv9c4DNK285/fBiJunbTThEiEc5AB7x/yVX
A787pgDvA/KpB5IBf/1st2a+K7Ar8VRUQf1baKbnmrE8Zhv/SOeO6jJ2eSk2gA4wp5c9eKitKdjR
bFprOZEVLjRq6ipfueTRTNG5CogBi7s8aG7ICEzO9NGdXvAKu3CaqSeakpmxNcBhzs8YLJpZwczH
mlp76n3qBGt0QCghkFBFBK0c57+SKxrA4N2aFr6vtsXqL84VMI5SdaK3azSPwV6tUu8w5Z/X013W
hATBRGIZJOBgq2rXZYStZe7eLiJNXfR9vljTfaVAG2iVez6ZRZcxwtiij6PR1wIB2B7oEId9FXle
GPn1IpIS4ifauYaGfFlG96MW0Uqmrs0qcRoDFuDsY+cKkZX0E58QqmqVykd2FYSZBtrrxvipLxIq
IGC7xsEVnnIq1F/fNf9rMU09qGkTSll1P1quA8PufjNQQf67apTYl8JY4scLZpgoa5nX4DYbLzul
bbDaTKuJbTMaKOJLUa6P4EVWkTYtrdWBTmvSGej7jJfAU/Zx44uTdYJG0K1oOJZKd3l8Lsmdko7A
L3m59rwCgoPYwrENHF8eXE6Z4ecewPo+x7znbyfcCHCy4ld4keH9N9+Tn4V9/6WrYoUmA9wvkVeM
vSBHVFdcSwH+vhRDrX6Z3Rpj6qtfXypEWnnCj3kyQ7xn24LkFCt55758XwhDKhcT4junFRpm7x0c
S+yhSUJ2g5b2ya5BSr857puydIG+KouX/4zynhrx4FEIT2yfjLjHOHmE0oCAkEx2VHbi1nGUu+6k
gAAxyNZJw2ruSmTXLZq4u5gF6Ei8UrcqYmJLW6dLkQzeAMyjbemZo+GY0cMiSmhfD+nqP8886soq
sgbEEuel/nNu7wSYnxmicLwqHacONETldma2MARkbnQ2u1CSo9IhHHmSww0qIoTFLqhW/pYIjij2
/k6S4vIm/m5t9LCaROXVAjmuEKa2a0ZwReOeICJyKarrhLGUgVCdTugTYTZTzI70Q5nVe6kcsVpS
wETOChKc1XU/W131/Z3cyL/ODyeKe3mCANcp7KGEXwdmyHg6nVZb7lcn+hicMTXWaAJKJtcpbNEB
dxjQGEXo/JmD9mT6KsjgZg0pvFhZ1vWBW1/UgLepCYqesX4vUkBcf1tf5NxzQP78OvEz7qQFreBG
jXojIKzV3XZFKJP9k7ODYJnRhlSBWTfc/vqAcycRU36ebh6htQIpFtSXufeX05GYT030bkyZuRJt
tdtOFpAZZCOQWEz2uvinMLwr+Ow8R5GqO6H9yHZzPJW6TwCBe1LrpBxW5YWAKLwjMZ9KG6QmJP5h
RhTAtVHGJexCL0liaMY0619TnIMl6HBUlRMMqZvrtmdjMs6mPDLBrr0tJdnFfpHh63lvUug1s6eD
6j1SZychMQ4ItJwrqqZt1Z7i8WM+iN3AwsvtywI/y5rUgJTZg++2U4TaXn+dEYHKRCIBVce1ouWy
Sglf73oGCW/LTJJy2EQaBEz1Rp/KkCZovpOVfJuO79Ms/MkhCV26tBSbz3VQGlCLlrjh0cea0XHD
h251jYrbxepP8HRiJU8BWVtgDLU8pK57Fjk6ID3R+djdfSBY/yTaFFq8/jvk58GEg7LtYmK5P1WT
Rnp9h8A6d4tnZYIE+R5Q3N4I9AFVtJnxuBnQ9IQqec6SQjPbMK6LPzDV3ZimhR64P7n/Ylfo6ggK
B1T6r8BsBlzlmqayaKCmjjSoEgplFSvHlUHrCqiWpan3N7NSToVZ6/k8GW2Y3qKSqmKfDP3gHEMU
RsRhtOTbU1xv1ExrW20kcI1ZVHf4unCg+4Rx0OF6ZfHNh1GL8Iahk+zN72J0r3wDlsj8kRc3odOm
yHfFWkUPPSYteZ38ESY5n3ERz9BOcYUoRABWhb/R/v1kmbjSiWeQ5/Bed4Gqzvv4FnsQdPihjjPN
N9/4fGiaWM111wQxXaepwWqIPjhShqR1iSeA4BK+4KdPtzQzHT8n/igyIN0fWPUl1mlti92JVytP
R9psIB1Kf13ADMiRoblG7zFTxZQsBM/gKEguaYhGYnnDQmKIV6gEt2yyqCEMsE82o5MBUBzXMeTU
MmNI059lqbrPg154CGtdKTRqJI9oHNKDfNPLZ2TaQGeqnDJWmgs2iBvWFI9QrOetMewHpQn5zhPS
K2OGePMDBZskn+muRTBu+vKSz54UBE57GN1tL3pJrFYsDxvBGeNZ5AicMOqWexWojBgKof20yiFf
jtvFH8P9Esc1WG0lRRK05yGXk/i/RtELECVxzmPI3xpK7qz4MHRZU9NR5RRXiBnVh/cOo6JYZeuN
xB9B/XV7+7oBHI56S7M1ykZpJevk9EeevhmD8Dwz3yThTsaxbHVqyYDAmi21fjkuDOK8Rkypn9hh
j2zWAJrOCaeN2fSfjmR7SrNUc1uyDvoTrBhr3zf0I68pR8GhMAB62WtIc09PgyIRQ14thaLl4FT0
tC+qwsd7MCLnJT48jpMK//BpfsxMIYArnNWwpG6olOdNfSWFjvlrUAuRpWDXd86N8W2Z7/vdKogg
IDiMkg1zh1upF3vGSehkjOAPBlbt+Iz+xUU9AyfLJ2LcXMefDvYVPKsxSCH5ees/tTPGEzpPxxF/
XCptIClr3UHrRW2qVGAuYG96++PLZLqSbpRV0RpeoiCHkqFFJ7p8IRk/xkSVAppO/ZjgzZhri6qP
0w+h2pXkJmhGDBXNeG5T98dUOkJYZmT8SG2Osg/8guHC38Pq74h3L48XU0SC3Uywiu7V56Cv/tEP
eys0mCxPDpEq2MNFTL1XCc1V21c20iEDib1zHtz1bVOzSRau2gDdnH6hKLQBHIu/HJStkInDPKuZ
tyYdITIoCu8CugL9+/bkH94Zc/cJMsLtDaE7zJm7w2hCkLYoEiFJ8yiNhVK3qC+X9cS1P4S7e1vr
arSZ6vUTvFFiPKow6DKctauMnzoMyrTXZnJf9I2dVt+aPWJeQkhekAP7ightODHfRml6mxUI2d9K
6TJcReNV/NLhHU+DUU2Xonoi/AflfnhvzF6PIb7JhMirVSgf1mYAIxE0K/Cpe9Lu7LEUHoch0p+I
ytCA2AlwKBYrzUgFwxrOHRxxYog4g97nOFwNL4CmOJlAq4i5vo8Os1Fsu6eI/qEhnYTti8mQFHSl
noxz02gKfk0cgHyJtUKsHLbcjfMGIGgMs3nxOaNJW8/Pdi30wha884mwadXQR7Ty2RW/bH5ewvJ3
vUSNE9zg3J0+hFYBCSV2t6uodAaNZKKRdLBXQH8lQ35nPX9nQDJSlUt27+U6du5ySeTg+Q9DBz8f
bENE5R3iVIHaYzRjSt8mPEwRTWDfPVzdYM0dNg6lmmFTHwDDPagUQ4GitWbCurOes/68EZ9b6Fs5
v7V7m+luWoL/yu8iO9Ha/33x1vwdlhyes6oD1Y6LoZMEqdVttvopvpqBDXT+XQP1wcCUUieg5xqW
NnwTVwyXZbIqbNiYeSmriws9Ba94mBIORZENQZuoeiqH61+nHaKndcnFZoEuq3t9i/PBMO+VnTme
BZb0Xf4tF9YfvnpaxciqaWBKyX+fkrfDpJhr9BjC1xnRRnQVW9BDdIhAAch8Z7VoiUoUvJSLWLOw
iGbkZBn1AIN6hA/Sf92UT0QXuSL2ZMuJ4JjxsxCHpPKhN7LQKt2t0H5ZgkTgmRBFDbc6RroOJe/J
I7cZH8AxFPU3atlFoeCdQyhbuTlUaGrpObU7KLTJzoEhwPWl1zc9BBiM1mPLxb+2EwN4BqVuqakW
xqGMvfX2GDN5B1KbX7Zr3Ue/ZrXXJNjr8cm9etzOvmPWd/QW7f+Ak73FUOxcTM43PQpW3esc2NXy
64oW72629jrJ9v/maYVlMcvCPzriRDjryAj5HCOgSM5gcEoSQzcXNgev9/u5Ikkwg8WM/BJdvBbn
n39l3XfrdZFFOckbN7TxGhbHgNjGHpiUM4Ggxd77mj+1DwlzaBKMTvx3b7QMBGyqv2f35YUA0VSr
I01GJHkVHVoy/FyFGQgdXHglNr6nk+vUFND6nF5cKZvx/iGaufNzKS8zP0FPBfY+RW9y28gmIS2l
//PCwjq7h8Ig7f/SXA9tO39+2zH9Sq0HbKpJOmpl2FamGLsBsawdzZAsnZPw4zpVWDC7+NkTwiYg
zAlTH6gQK/E/u+pE8f9DMCKuiftZXN94Iyn6eeNJALHXNr9pb5Q1fDFFwkxrPHaPXMg5Bd+Cdp3l
wFcJ/d+jpgg/Lt29ERVKemElMc385wiKJp8BYZkJoaoThIdI8QptesIMOyFZL7FdcNL1k6yypbS2
Uu740YTheJ3pmfDTftvfgGZFxKArTWIy8HMYEYKFnvRRKyPAPtyylLajKm8NozEguuD+MoWzy0Nr
TjgPRQiYSrTTT73I0wWDRSHoiqYKOneeu3b/MWkHkxagpB9WjanyBl7bgFt6dWWALs8X0n8585je
OBcNgO6mzfhAq9jz5UZ0KbAmH1gYRYsejvJANt8eVqmoK9QCBucbw6immlo9FttsmpK//C5have3
LrQLQPv76gDfupLLYayFJYGlWgoR5QxoHDm3sCtRHpQc7vPYTpH2xcabfFErYnxA8M2pdD5Hni40
bv7dsz3UpHfcQ/iD+Fm+TSnYN+qRop5WBrhh0sso5S2eNpOT4PFWC4G8XP9E6SU3sf87JbBLYVgH
0ILFQbkcd9Z+s96YNe55CqhPAnPKz1duNj8tUxTuPSv+Q0R6aym03DistIcJ4IjNF3bmZipKgW+U
IrarM8HkrkXRjiftG7gcI7vvNV0LoL++jTAEgTinpzfsiXF875L+Fyxk0s1KYCASjk1DigT50fFF
aR4oYx2OKXqo1CNoDEufflrIM/msDAzfPeAaYHXYFMBcl560oWoc2lq2nfjhVGR5mTYUSCDT4An2
12RsxvCR4HSjWMUT/Zd9LfFTCVCFZYpaYEx4MmzaRdMn7qIFVoJVAcCxxBVPIZI+hGv+bn0yzqIR
uuIXAYKBhacGaY8eOYFOP0koH9fpCH6bL0RYd5CiDNCUlh8cNlFcwZxLT6hSaJmEIIkJSQnVqpQt
lUy6Q2+z34kULT3isiEpZ153I4m/hn1aDaGv9DFXzztqk/if5lOHcRuDyxkM2sGMAZLAOagpgyJZ
dzCP86Hb92BMYVUpWO8yYfctI2muZpeywxA9Jy8YbRQAGPg+o3+E8k6yZ76hfZtGSPVsko0tG4jw
lT/AZ5uzQjpIvTzlZ5s2MIA0REZnLkCOfxLsx/FAAb/MbLQHvTKnyod1dK63WddwvU2qRPrE5iPB
Xv10UiPrpcvkrU4HnWsE1WE2LQWhDef3eGiTZ9kGLxKPB7u9kyAmn78zS8fXwcEpVfX7sb6h+pud
egUe6pF6C6kiCQoU9UeHZCL+nJN3zApyJM0Aa4Vfkxu0WXGCgTwueFsTnDjJqZxzi/Xz9MoBsdB+
IW9EaLTtoMCUJ75XJKT46C59nWhw5RRYYODR3jruTsLevccdR4luX6zA7febzbNw2z0KGu1r+J6x
VaQi+ZwSjsmFWWC/CrOyWB0Jh24B01hd+sEr6CqQNe4pjLH6DDi2ts6rcwVXMlyhUvxhO9dtey5V
i3Cc2SBrXGJci2sFvvIy3r4fyZbgyriD7yXpXf2PDkiMoC6J4w1bN3yNsT1LlGMhBGZ0ywSa1D9S
mdtumJ2BZF7SSAI0cKx+sES/ckW0HkGu3hvtMf/ktT78ymqKw94mIJcK21Mik5kwoe4tKqWEA3/V
6BT9FINpJDoKHgpPbNLHuOAcujZcWotYrinTD0to3iQGVrHCZGtT+ZP+9mPRZGs75fr6rQjo1ZfB
+yVAVkbueIeSPLVlxPb2jGlYOLw2gS3oCfKPG9OoLgGujHEpN34TogqSpybyGqihD36cbdv4p/Cu
GAjjfibj83uOQMAo+VPWgde7Sqmav9xHTFdaMACemRhNUwNz0xZuZAmy/YcXm3fsbJlEBKnTTkLh
OjjlsCnDVJAWA48qgXUmz7uDxxYwQlxKINHno3/8oYEtffv6YGQmzRh9dvM2KPeyxzDjwBMJZXk9
OrO3JbAAyzT4k9YCJUxI9zpSCMT/J4CJiRurK54/0AQCu8JMnZvMm7LjLuYuM1GoYg71xjNPEYVe
/INiTVNe5EgIDN8R2ARuE00D62DI796LJkh0+L6lXH9rAILLD8qQPW6OneACBtqeSd5IiPBwoItG
kSVbcXQivWX5sreMg/JYU1pYFe/U6NizdFlw327bFyN245n2ZgwNh7BtRa/0MgVfZu4zXw7F2fy1
BYp6LhuYEA/XiAqBoNbeu4z/VMma5n+ufkycmNmrCyrUk6eEdbA41Z8CifTCPVhD1g3yaSVsEboO
IT92CVpg6ChhhSyyWT9mExs27+uVym0MQETiORBoRJBzJatt5M4ERBqBWtTGOaUpp9b1TyEulDRn
SKEwjwB1lN26apUDE2KrlndCcH5SpUpLFrbhQhPAI9gNgSK46jLWeUY8/zhwxcLVakLqbDstHwas
tQl2axuTCT0oHD+6z8uydVT2HOiyi2O58nE0eIwXyIpmeNMsPQu6RlgpVKgdw7kpt3fQ6zZE34jb
WzFMCCbeyCg8rIkH7XuAFHjehpoRNLT0n1dQigTAumWmBx/mx5AvJmnEGjRiWpGBavGolZ/hOhHn
zSH2So49m7gHj8Szl88qSJwllRhAXwXJAjocH+k17VZEM0l0vDhphMolV3vQ1Ew64XekrOdIRj7t
sk8N3qLtTJoePwEA0kJP/32+nSITZv8wRZAxF+CXYnbM8WEvOICBOK6HyOMxvfINNNrcHJh13X0i
1fCT3kVWkUdc/fukTvoBxUAEkpaB6tLcMO9hn0suAMHJkPWsZ4FdHByo14x2+lAFks5AtlyVXQZK
Qu1k98RN5vT9h72GDYc/7+gK4/vgnrsL74ksqqjLq0w34eCSII4yWBs0N+JcUsVX0YlcZLVNtV4Y
b5X/bEvdkmqcjPfb+SU2kht3d3DiYff+VApAFqiR5QwKx7IDHhi9FO5RHD1WWMNHwETswunlhptp
0D4VXvMVSLQKFg3jZpNyMr3jdpyO/csSSqG7DV5be7pZJWgAwhyXsnuSu4jOCjeFYl0eMdodGGel
Dar16iCv1pTuCM1OW8yFJJaz0jVUh3g+iymSsFX+R+tCF2s1JQlOl1cH+2qlmkX3g1dLs+5fkZ6P
sP9wzSvtq1lp7hx3tG7x62CFiguVgen6eLwJFSYiIF9XT9V6BPV3oqIj9BYFByRga7FXCiHj4+8V
BjUVTJfu7Zsa+IHZJn5UsHOGh7STjBa/4DjSyifoBmLCsM2iwJfG0ZjPS2hQcaHPV7L2ttso5i6Q
rFLnyHYrOzcD8pQ82Hk5PmmSmrSdASRV9wY53iyCrs5haMxNsx2r4QtKvvUDthBhY3c4Nwz/E/Ts
eYri8ZW+jlgBEyibA4tOI+5BNOXl6S1NcWYLhlzL9C/gUcDD7xuVXxLOvtKB0q36EZ8M9Zli0B8k
PTyLka8kGdyvpBS8qagxESGuJXArWIDTh1ew6FjfpsqwBurGSCmhtTb+OtBrogDc8YNLfaMWp0mf
VBhzTUXz05yPcBc3p8A+8lw42s2dMvC2LZ1PmCApJfZm8rMKveULN7j5e1YeZd8VUy+tkjbG6IJn
LVOhk7Jf1Zl5+d627Qy0oc/alTT8rEyC2i3qSzNyaWJIwTQsBBG0Dx3B6xrNzUp88+czsMlHUoCE
+6nqFknQQAHRP5O/17Wsi5dMrk9HcE8A6RFUW/nNh93AbDrxTNotFTwadZo68Z8laJJeoNFUcphu
8aAL0M2bdMHldMCmVhSL9KIFsyN7vhJGsFif6cAyNurCa4uBnqogZ9YxT7kNrFJf/CsgYQ1dNhaH
R61ol8maUz2tl9YBy5WrKLpV7NF0i9LT2ThO6GjRsVEROKlSZIWb4s5uhcUTJSSj6VYFpLEE+lMl
BrYIlrSjVx3hHwCMJGn1xiLFoZrNWcBaGr6FyCCj9BQ3T/Ixop9LZ5XlxTxHglWzoR8Mc8mUOiDw
svxfYwY1yitX7oKXQx3Co7TdkplLnY6I/6KE1BPT8nnFkQR+iPBeLznZrzx5rPaFRKz0IVAAjlCY
DN80EGmYeLudr4Qylu8381k1w4SavM6Hg5k3R4NRuLHr2v1AQWDTmlRffQGnEBaLxkM9KQL94BH3
DSpwmG0XMvskJHp5kPZMa2TqUUo91+tNx3z78IM+JRDVD4CAxvbzcy7UiagyY1Ojnd26QukZ/yQ/
fjTgWwQlwfP18ATHz57OzwJH+FcUeXeK8iIUrGYAz4wz6IFsgRxtvXaKYsvxkyoQqMt9lLHSlTV2
KOYFBjq8pEeZjhBSN91O4miSnIqF1CHCj5H0NY2CL25OscH3OrQUuEUYZGnfoOe/tebEOITpFCbd
36jrawj72uViS3U1ZtQSyjgfCaguyf3pX/y7nIpvimYiGlwsGdijpMANx/J3WE4L8zxwMntRv15X
zOhweF/5wpB+5vYvyrz1OpXvx2EBaU7a05nutRIIEhjSIobragxUr2qbhXTpsC/ts2Eq6CRTJCLN
aSLWxPrDlFNQRBhQbz6TsqMDSQw6s3L8yIITb+HEe0w9p86cUc6npxm/uXZDGaRRDdPMfcmwd/04
arR/vXxfgQb+ps3U/ggJAB5iUiKcRqtFBeMj/+9tT9QcN5K4IzhGG+Sg8ysrFqq70M4LVaK2neRX
cjid10F86SjomNvJF+gQPSHUsDcC60HxtIgeajF8LkYQGXBY7U1R38aGyfTEYgTHFBA+LmCdU6yV
3cDNnMulcjvjBxgJXFr927omQEQz0Nztl7nYFdWFELYvEHcF8j0+ULLuDZvzwHQ6RrlYWFlYw5GZ
f2yqhWzNLyek4z9+E0btBUUFmIP7Q8gSUAl6h6rPMCKR1kblA/KjQ/xJS9ZxIRzq5K0/UMovxTqu
gSRdaZhN3nuaRyiK5MzmXUlpcQ+kwWfnNdau2QWGXmK1T5pTWCN1X14cR7Gm2uk7FPYZZ6pmuQ04
8K2yXl1XcGyN2S1ODSFV1e2SkvdgljOPHRKSE+BV01GdGwrm8WMv9B193G4j9c9Fz/HD2XLVMtl5
dDHcS+w55j5R+nJR0DXlnt+i+IqR69VC2pWYIquQ5xqjPVp3lSWR9K5UtQLl13uc4Lfe1A0vRAtP
8LEFcldE1QLDCeWkJkzWPElW1nAU4WIVZGmWFwdxlo+MForyp8A5Q6u9L23gCUXZXThYoFtHDOwX
rRh3cnz6vpr+yAvVl/kbVM6nnlqX5HA7Z2qDYgNJtnYTlcXIwt0JjCX1wMvANX3SHDyNWp4B19V2
4A4fXTEHJ+r03A9RJOBvVbtLJG7OyEVeEo52SRaG4iK42ODe1a9mnvYlTlukVzyKHBmocbXIY3Pm
8OLqyKPXacAoAMntiTlN3TzURzXtGWPoiFUxgAXvrAdX0/76zuNWGpz9VCJOH65PzGoasmLOO8tu
LqRPcXUAM6BTu+9QyF9e0nOQ1iaBozFHoMYGCFbWgBGs3GIz084Bclr0ngUQR17ixVOCXOdok+u+
LHSf1WknPpjw3YV8+sE/AANjOPRZ+DEo4dRJj8imsSPrcbc91oJKWTiULYEgSXKXBPzkfLtj6VbJ
Oh8ploBZG3zVRq9y6ZmTxIGKfr9cYwPVrIE6gzw9PxXEx7AozlLwFr7D2nJuGoDKq+XyHVDrUlJ0
ZdPKJFXH9sIa3BAg71PdpBZZWkSa5F0sAW7/k6kTwP0G1J/L4z8E7B4FZzl3D3AQ1ugFTUcDC02S
Ht5FErz41VBe51WcPg3lZiZuJWa02b+HRBiJbHXDDp7JJzTpDG3xScSHYmToOMtkZdfZHAY4/QCg
wsfuOpg6EIxcLMU1K5Dg1Ga8NjiVqtfBFTucelrg9u/chUWyBVmcKHrxNR1svBSi5lJk/JG5MfbX
73mRv6DZCphlwTt0VqW1kKILTRZVdYgKgLiHfjFnIUaf/zQBeKw5Tn7y+tN4bA8k9uC3h67tZcmI
6koZG5KZPIuLJZxQn+OzfJaU66hXZsSS34gnWK5AhMpY5VMcZNfUL15eIRbMKac0DBKE+S0xUhO1
etJS1hvocfJzy7B2ihtuQXucL6OkkUx5npD4Nf3c6Z1wYTGlTR6K0M56Vc8txRDQe1n9Fw5h49k6
0eTZZ+p6dTdzkQLmRpVLDglllOllxM1Di8IchqsaCXC0owrvsTcV2KtzgSHH6kHAzfyfvUnl+XwA
SNluWKFGUOdnUDK0ppqvZbeQtEOgCiNvSqPAiRS+LNLDMoPKpAJ4HN7Y35GaouNR5aI5+2eaGUix
mN1Bxdls3XKdHUREvF0n/caKZjdLWWT655MsTLbPyjjEBnFYFEFvAON+lW0WN08MpzFfnQV2J0hd
Jk8t4cTkxe/jD9jpBiFMOzIA4HwksRWl4ZmNMNwY6eIbW9s0HNTJb39J0LeuJflzrmOg2Cf1Oh/K
A1VLnBLVzxRUl1/qpBC2E/zXjfdLrUW1BK+M2BlBpHO74G3NmLhOHBdFgnftSil2OkM3mZxMosc+
BN2bEl/5hIxhETMqLTre4FHtjosx3fF5SoPLgezXf7laAvG73thGPsJB+TTyvR78BIhtyKPrt5zx
5dvBhe/CrWgmjQj4T0gm/F1AvaKpK8MJbPbe5vFXga0VbGr2i5Zpv+AqSj3AoE3zx9oLzOOSHxb8
q7/fRkr4HtXal3yex0UcBXYyKhmgYMx8gFqElwsRKPJSuwCu5JW6qnNG/xhplvd5bCOvuPLzG6Lu
//z2yuy9hk5i/jfZ9DczNQynG3pd3qS4hbGfnqwmwI10xF7KE1SnDXKfJfh4yUX9ifYxW3SnITS0
ALPX8eqLYX7fweFw5dsjn4AINh0rBSDWFTZJWrBc+4SdFzCtAdCKoAAJHa0GwjXTuiVHAHI3+RQ3
IG+Uuw+hP4f6FdP298WpPeRNJ+sD7+6rE5ez5o4sDjcUVvLG4ImN6RwDXakazFJxr/j9lnu+dGMz
LMGceOt1P+V9HRYmWqQxa/ipDLo8jruUB6lxbFktL+7p3j0BEr9VzvWLA2/eAUWpdt/x43sZgQjQ
e5wRImUiLb8zunBNFlVVEABdoBu965lso8AazQBpOceQZaHaMgHnzfjyEmD7mfqkmClnOSSWmn+4
MyJN3/fH/KEKBjhQZbqzCCz/vgCUVu7MQvSkZn+PGMMPGPm+d5Wi3pa9Djqg2lFA3PQyWjt6rKaG
vbrb5CfoD/CWjwGg8j4q8E71K3pORmTQWR49fQ5NCO42XCRL1bw19jvte3mPHzwL2qK0AZtlDikQ
hUaYOddtO0HqXdURJ9mPeRADxFoTsE9p2vG6fSCoNL/mDL6wxl0sCjRxPrJrF7NVeKpuwy4RlhxW
Qwx0wniNn/sd7RH+dqU8S7+qY7nGQYOMGI571BbWpwZm2GHJf0+rSeMBJ+tR1MXYKVFO41CaPklz
Vk2DIkEaq8HmBMqT5DlBfjgBwRE0cKaYwouJt3/aJfzgRCTCtvB2iwTql1benzdul+JDPnS4YjrV
Y9nBOsuvK9AlzH6B6aYeAv9CSM8yzXnFAt/o3U+mjNR4dERZi4yb4erWpqq4xSJsiYvlMzAl2SaE
WJOJDHSBk4qBQO+p0GXJYs59p9S0wmB2gXT/yi/w/3rv7vxq98cTzDD+pLC5PHIFVPhtxDc1Q3nN
Hz611QqJAk7B30d7ObTT8qo9wt65phyWUY+ea647U1JhWH0sTR58f23jWdcbVizlPJUjb4QWUB09
qDYagIoc3YAtM9E55BCYtnvoa6eeZUM/FZMSsLFlYvgfO0P9+SZEbhq4LdiP3HXKooCrLQdeqpLa
o7TElDHQoNon7zJzqngxq0GSZRPO48NSaM5VU7qeyIEA2ZNt8i+hiUiZDSudeixvOZGB2ZgsKIrs
IhCD19hhEFFh96Cj4+JTxm4vXeYzNV8u7lbN0GHd9kOMzEe6CoqoQo54dcNVCa1kEuZ8cO3dESOq
bi5MPORyVcEwRvMmhGiHyZA6I95+7S0/wKA50X2qRiqsrYkLLmoSoRiEpaurzS9YUQi2TOrWoCSr
yRXKw24HsVbUCE7Be/VI6Bzf5OxRtW8cFrYwMVzV0OBfBcqjfGoaFOzexf479KQ9MiPklL/kz6zY
qBdw2pG1dxnFQ63TU+7p6IE09mDnWKsqse9c1AP0Da11oJXEpHQPC5pADQ8p5vfSZ7snLpH+LXGF
hroLM8x5Xk802ccgAc8QqdUeDLpibPnzAuRbwCBFIVIuTvE48iNnRFtaI6CXzcSmHX1Kkk6ACyLt
BdCV6o7DLKxHRewh4mtt2SkHYxOmqfDN5TjuIseRC/Ks8rXVO2WY5NlZVYJATc2c3QaM5gNH4c+R
w0UQZ6jTlzGsI3lPvfakAkcjxBlcJW7VpvEk2uBvzFgMhYiubZCHq/VzkqsPf8EOtpLIT+vGWrw2
2P5wjI2oEiw633FFAVus8O3pB42IxFc+4VijLO91Id/6o/QAdYjUT0BiDV1Fw3Q60fHlPJwGEd8a
uVP0QWTVMd2WWnLCfOojDPpD8brPD7pQIQ4q6kCf9k+3v3IlZ+yEppuIEOF3VXYt/+vkwqZEthNi
FaH6elVst99prUUtieOSPv0oqXz5YPlZtY1cgrCaUMFILHNgFeweHlD2ufhnog0lBAAOvTjtqCIn
g5QB3MgUgUNiWaUJdzDj2p/DCZzME2jhli5tDe3gPSulJhWvtfcZcU8UNjHVrYxoAlCk9zFXgWRB
Cqzj7P4L8gOiHRTO/g4YH+pKqeac9ctzzU5GyEbOhZGzIiyh32InFzVkGNegYRPfIqqNzFQT3KHg
Us3xNjiwgV0+x98p/kOvZZRx0oa6wmYUxgqWh+v2661vqhiyWvJ/V7c8pbJstFSzb0P+Yd7Brois
WGBcOLBCLjD70WqN7VokOPpgktXIy523GE+56VFMcHHCLQrgmX/xs0fi8SHmuvonytotFJV2IJ55
z4K++iIQc4VBYPyKmxC80Ybvk5xMTjAxf5lHKVk5YiA0+lqd6BpehSfkz96OGXPPsnSUI9Ebjh+A
Fk8IVd63oTMHstujcerAWQjWKwLMNSf75ED1Zfkxt4G4jLBtetj+CeWg/PUD1UwDk5CZ7bdY/iSM
qW3y9/tLXTy6B8h5HvQKZ5/s7IOD7rzJmYdhTJak6cTqdUXoCTBb4+ompoySwSMtEdv8ncVlNrry
8A6uOEGJ4zCBzf8eP1rSyzc4ThBxL6rQP+6fD5eqXpASgQgBLCkHgyiOJ5CRVile/na3ktuHx1HR
cYrNlBJopwXz33Er8m1HW+UnyI6GTvL6v3s58eIDG2UPD9BHIhF0Yw/azCtgzA7N3GB/ualMWrjO
kh7zUraNgZbjo65wPjlb6i8jgzytiUxGOZGqhF0KifzvB9AC54aS0DUuAFrCkDY+MBjLsKy5Qcxq
1kENaGfZjwng7jmvkIGKs0Hc6r+ZT1wfsYL6XjMyb/EKC7/UwWdlkho5FWx2LqG0gfQ2/rHJdR9+
MWmB6rkNAVgLl2Imbhn7QJvhqw6C/Y6eDRryf039K0uxIsXBYzSQRCQj3Rm0JeC1vdLBjWcvMJR5
MbOSzzDL7qKxkGYZKDWHPFh5NT3c87xo3TnwTvCj2ogQNs5lqnStltqgF5IzmpIVdWDsAzGjg34n
RDLsfNb1UNFAmE/I7nCPDRLpN5VbbWHo0psuZIKHeWzN8LukEiP9QDh46cT+gz/luqDrw0Ra8gUI
NP9qMFL6xRgPC0GKStq6N5W5bA9HvzWZCrPrrSHUT5X9OtUWS8XJ3LJeSMppqzE/Tg5qYkQalJXM
1yZHCni335mEgubS2u89RFBg2NJ0MWRppXmKxEVCD5o+iRMMu9hIb3My2R6OVm/pDAFssFo75TVF
EWdawVQYjopxIR+RmOIxHa+kXrBmx790OT68Ms5razarsbQ8U+BVqfsFeW7IJJ4qJ6cOwMqsg21M
0sJqtK8aWccgNEVZLaWms14qKMw+pova4+J9fNBIVEbOZWKUQIVkdi0MmozgxNA+Y6T2Lfxq53pd
PIkSIdM1KysPTedibTbKt1O+o9dQWkdBoILD8jOaLI4VvMu9/rC/2XZnmgVM4XBaK2fIqSyUwxQO
GML+5mrLDLbarzPzdyqg/naFkpPvSk02fpo8stai9XeRy3NgWcKPy4cTEZ7KUtTLuvBXxOYJ0q3A
dPh32BwN5pPFX70qhNIvHVflp6Sucao6BYDaEYBibQz8cQ3mV6/815XNVZ5ZbzEJZgu8FnUERlKf
bZWnZBcLLG1JP+WUOh4tEJCzHi2pUwhn8wiTo9sQUBiDcRW2zpu8gHWNxoIiWuZmGoCmB/IiJOgD
52HnJxZy0UDyTSyVPz160MJ0oJQ4VGuVQCC+t2pOutR94dGLaj0jer1YkNgYq3gjwDINxnQIz9/H
ko7bx4zxHIToIpVlMGgYHPHTFdpqPJpfkEBVgku97OA6RI2LRrGuxy1+SqvzEuPVnIKLCAQbD04m
G0SkVDTcSo8K1l00UM7mwOZXBeviSfh2z7iX0jFfb3Bns3thAZg61CKVODVLX/UEfAKPPmBINuuE
sAMKlyDXCQOrGFFLJ0AYeOdS+TwY4LI8n/NlCU6WJvyKDrQjVRbq5FxpVfHRFA==
`protect end_protected
