`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B9EdoYjgQSD9gDMqVua2zJVflRHus/LVjvgqriMNBVhHK/84/U2ioEKVQOwfFeXzEQ+lX+hFCLqk
IZ7jFFR3eg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RhpaDjajcReMSslu2NKOwc2kbW/sae+dRFDHfVBTDCkPzbh3mSiP7TZOBqhKDGqTB6232MKVx7qP
ZBtzaagM5AWVdbRcklCBM/Kdvk2QRYet2hF/9C2MMh5T893aaMICNr83Nm8Vp+EZuwMrlQi9gn4g
ywBMUWKYky2UWYxF3K4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EMspBr3PE9iUGaTBx7AjQJAXSHmvP3RUIoqkvAbDE+yVNcZvKmwd5igMnbjWzn6mF2c0q5bTEPiV
SW2sgdg6e+BWLSQSGz4p9DMI+GfIfZaVwwQEDESBje7X4DTUoGoCTuJszgnSgaxHrTunK6Mskti9
6KrQ+39Cj86aIm/Se8nuNq0dyvAGREfF8mO1NUC0gTq7uy5v/YguCmfE/DQabE0hSg1HMsyBV/Es
GiQUjqTbeVVWXfqfBUzosAXVQKO0zqx58iAqNL7CvcGEpsb03lni7FDq7sA6yXUkDI0QOTEsrc65
s6ZtU7tJTAb29hQhoHqIjiGrJFezQoQSsaoiug==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b93sxpNwCcwf4KNpCEGGFkec9bpq/IxvjyBQsUyVkA9gs5+mZCPe1ZsIgPAcV3LuAs/hO5uF5ZZg
8XlLtMGUzLOqudI5PSmMsrYFDtN3zZH6HVVdrqx1SI+iWh7n9QVxAWi0Gb+MTGVlekns5jXfAoVc
3u3FT2heMRrTJpych9M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bXZyR3Gjk3qu1g2YuorAQnE8wshy1nalVGdBpmgUZ44y9It3o4HVFeQyueq4jESAF2Ey1VYIbvPD
74ozsPhX0ixRYVusT9MV8PD3YG6LdUBXI17bxA0LAUmItJloxWSXa+t223FfWE7eNn3+E2em1yes
DofEMqIUoCSM1VrQfdWQHWipV5VENa16uK/O6WvUpm9HCeZutIr06Cd4/jMLDVN4zK+BRg6PzYin
7YtmQvIO/IfyaTOOFuJMXbkqdaYK3LMmByLBTTcc+Ph+MSoPOSUz0iJ+rEyUD+vUc++9MXYxYO1R
d+2oGZu//gKeC/sSjsNzj/WkgVmTtfVW9cP/BA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AskrFrWXFM7AzCqlwzwplr3AKnGiwwGzSK4bMSSxCba2xMWeQ3z633VSAcApQXs38MGCxBDDSYbX
nUzKzPFlZpAxD4jtBhFZhYrE2rfiXck3GhW3dp69xEgpUQlfw8i4t1/+iPNzpGa99NBOV/7wTUca
GQByFwIqxvt3bKLQVKoSCzYzVgdmM4ESHX39oRKLp1CBheiJrFmXRi0x2ea1efHoG3nUywaxhQeI
YzkcGouUEqPqhgI3U2ijlo/YVImbNvFBcG++cJWa4jTlqPyGPe3ENw0VgoihgHcOmdTWUcL0cLlB
R50AncMkumkCzB0MXaTqW4ee/PyvqhHRlRf5Bg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5120)
`protect data_block
FfpFEXU99vgoUXkUYb+7PHE2tvGpqRWuG3JwbFsocZV/YYzUQ2X6T2n2u+KcDaKlqjvviGs5nRI+
K5w52mS4Ac5AQn/Z7raiAzjfbZK45eHtR+2eKnEKqI8b6SktxZui+uszMKp/7shsBpajWlP24Sbe
XYlYNUxE3rYrCmwH4zghspV2N8DhXCRhcCemgpqeORg43+1EYERQJ9a1vqq82dL8uoloJcU00VO4
fe9teYnQ2efNjPtL/8QsiklonvBa+aBfsVm1G249Ow8x3jk8JZzGWd2HlZn8twTaly4AezVMLZg1
eU6ogMzgKRb+CDr5OAqfdDDKGDywIILpz/1+HzXQsYpzytwXFxWXIZxaV2/8sj5QLDJKvobj3zc5
dmv7eFaaoHSXg1XuLtIH2aZFxjCS9hUyktftt5MNrIiNDjmM/3sqOdRPfRnt7VPUvld09d8GNlMP
D08UcwmMgvvnS38GuoxhxqPRWugUR4ApK4yJrU7LIJ0RkE77qIu4/kTP174MfHuJkIv+3KWwvQVt
4x0i30iTFoaX8lxR9YlSQ0Ve1YbwFPA3z3/Lf/nvGM+zOq2o/ug3Wo3t4yU5pUsubAmdP5zGzG6y
MRDmG3PU90/iTCll4alkZqTunfMkFvFcPmSpRAP3IbMcwr5qTdNec/NePSL2DdgVkCQdk8aWsBRf
PJgLhGcUAib40FYbnL0vlFe6Q17C05QHzgjm9xRqrvDdannxedDWw2zZYm0gU/lmRTqLWfNqpnTK
R8vZk1h2fUqyvlkTIYC0PhKqEqVNdNBtWHBv9/h+xE+Rv6vHjaj0XyS8FVa2OdC7sg5//2wWWs+6
UyQ4UHx5XwnIO5dFfqc2wGwQ/AttO9QnklzpSbjfCjhbsa95kQowPGOGvDyn9HQEMQF66d6t8KxY
RuUxs/uMm8vZg9ab6tyLmaw2Y0WE7IhRye0QPwD7jfoV1V71goaQjg7Sgga3YC3c0qPsKIFtPwQ9
lqZsDHYWzaPcvPDEh9k4uFpr+6oYEpnXZRwwHc3J3iCcbWRtNK4S5aILTSFF3SH5k8VB6yyvzvLb
wcLUFABeK6eWVSl7qKTDDypaAEfUOpdp5LeeVh+Gr6xyzNdy2rqUSBw0PfB9dPCZusRGpo7tlUAd
/41Nr+gMNDrOCWbLpQjQALM1ZFzlek1VCW6k6eyrshTCAmEml/D88FNzdI66aECvTzhtr0Teu7m8
IQM4a96a+sQ68l2gtCMbR40WKYsdA5ZzYhP3PfpWKgsGI0clb+s8rDSrIXQ0jujNchxNkbl1bCgj
vmhp9okZ84hC3bPtDwLyE2Uv3KZMqonzi0YiJD0lnKqE688Du7z5XhYJiF0TetJEu6M4rMyl4S9a
H7gefztuIJARZUNMEPNeiJDclTmJ29n1xNbYvi3diL0xHCmAGAxfwgg8kXyOriXH1Qy6EAUHTKNb
/0IpmkzmU5ZE+/KN4RBxqpWdG15K6kgi04Cb93XZLcuvailUn8NbggzqYepUDxYyJuBTcnX+1D/Y
3GwfQz/XynGLlAqMK172QvttD34Q2lnSR35Gx1tLK49PmqlPSftWeauIFqxetam8+60gbdMc5Lc4
9nUXBzTJ3VLouVXohgVah8s4vinI0ZJuIVBml3SNlgqYOz61piSL5VRxuYTv1VzwS3KYWNIq/6xd
quKbnWzVhzmAych/uMRstnZ0whvDHg/Oqq+ecrgDhnSXR+tt/Bz1w2hNMuSwN5PmAC8lJcASQ/s8
arh7Y2n6AxCKzud/EbuIVI8BcKHkTIBUrsHH9haCVU6FRO9y2CMyvQZsvZ8Vkz3E9DNehKH1uCLH
0iypMxifu2BYS/9sqe/Zqkn+/R06uidTLI8rBA7qYfRxWO6662sPYYnTmlWru+wiVCqsNWPPZ8Ia
T3O3TmRx1rbwWBCzseVaeDuws1Wr3DWbh7MEOa4ACSBgwnmJPTiyvybco9TUbhDnp6BOy7Kh6Zhb
djrcKpEBQfndXMyuyaj1yg5NGsyM4AxTc0HPXg4MlE8ULZif8/kvyC7+BobgEiyV8p5Ru51PUTPC
JGfVoHBEAsSw5cBvgKCDX/kKhhS+J6/4VMhTJmeXuJ8xGanF88z2nPSsbKvJ9O5rfn9yKRDqRNug
NTyk79CG9hGiUkqupxhNLKoy0r9JHHNbjtut+zIwvdSQtPMJTG7KWnF68zcibcVmfLRToRsyNN29
r92R0m3gj2fL+/GuCrvLpEfhK8QQpHbieU+d0pL0igwcxmb6G77h3kUVlkFInJYplvUMvYTzZfdI
yVp8+e80x3RYxIsem0YXlp47vI1F+aLPxvRamvvDrwIJJ3ua5C1gpD6DwHJtG7gAcd6RBkpUa7fP
E0VXKK1kuLzRgjyUZj9URn3O0W5xGpbbHBoMHZ1bH03bKHtlHh8EstnSGjFFA7ZXqAOegCuhDQ/P
APNWU01OYdizRN312nHFJncVfM2LNTTCdSWD9UytEfiSyk7Jsp1qd5Xx/8tnsh567/JcNmZJ+Xpa
vpCgnI7kIO8KoJv+eH8/3B07tmWDgURTLk+U3UCM4QuX86cJd6IVNdOhFKKBwxaDpDrdFUICemX3
qsBjhbld8gTWyQxfbCvIONco1LdJSpOmpIpJ67o+MOPDJApiDLsPYygi2I+1r3/Qf3K76BWMUZ7V
FDCIPTPCIBu/O9K1hdRY2eGxDwXJKlGiKmP/YzQF9JCe17gBEtfqHuRrfi/YUGox3ZOevvSfQm6j
CYhhuXMfw8xXHbbMNrhrglxAK4E3GBNqlRQuzdKMzIk+cZUH4hJrdIhSliD6UukA3/c90si3GJ4e
xtukpLnoBLpExx8+0L4XAfXbFQyFbv4MmwDBPWzsFfzXhlM4oU2Cc7TYeRFn3oUqWq6W3wC7GntZ
5Kd3f9Oid1d6CZcfRdtNQFz0sy/kuHqJ5LQi8uDZUODCdbkCuOcZCX2IKE/MTkF3y8l8JCEr9leP
TYfCRBhARZL0Neo7S1S00vQF15QdhW/zP3Fl3hIAN8e0YlzIMrZd4IE4Epsad7EYeAUHdQq1J4A1
obrWGDsDC6UpigvYPqznGeya9kzAurcO+RfRfJO3IRa7/rx4xAiOkN6igWVDYr55U1T3PVUs0YIK
2pdLrTA45ihrwwoC1ol2mXwy8YrscxerS4iIA+N3simZDhoJbQdoPe3x0sAYmMnlFHdcJR+R0FGf
a05YY1/FR7nFUFWrZ8r59BV9zDuHx+gs/BBcn8gv3lQBKTL634aaJ1EO+buvvPpNpmrU2cNNVOX6
BvWsrymRGbWZHnks/mSys4fi0fTBsrLlGfGWqeQuO6WSh/U23q2tS/fG5Keaza2gHQ8F5tFjTJJk
s/ppl3BmFqq8IF8GoQbTVB4bPFNo+G3YlEm1XYRCPn70qgafdqrJq1Jg15kyJQh9neNGVL+lJm+V
xXG2VCc0UHknIy+dO3f6TBM8P8NGKPxn2tRH1DjkuNTVe2mQxQR2zRZOUdHLclUQGVQAEl7LasOd
VbNbFtvwxEZVoRfvehF1uz9OBHjY5ASoLCwjefiFmpoT7A1TsnA0KsDuPeG6B0ZyvQkenDe3/Kmo
5O/Xxpi5Qb68skmwaJL+HsPN2WrXBvlZXyLgoazipQrKzOO8VbEzK2C77fjaJY4wY0G2j9r1KwNO
iFqQW1k1kIjRPKQMqOFLLqtzU5wLukFBFSlgqED0kFjmFCCVt+B0L/LZM1/tcmO78vIZ185d0DMS
THXp+A54uUx7GU+oo1yRZndN1Wpr1M9peEeL487bGZmXHmyNbRyLSySZsgCTCrs/LhwvA2bga6WH
SmGO9FxbLFNiyS4xVcC/ubNeUe7o4BzKR8b7DIlHbi3KEd+TvWuQAuOMA3y7nwu7fTeKLB07t77e
hF860BFzVmaf+kBQnE3nib/xggl6oT0MCxsinQKv9Xx/uxuDFLimE82YMRQRtPAUoIGOsSswutTX
e3dH0VaM0RAfeIUhLlqnCT0OEjkPxiimNx9bvTzti2u+RCLgycHz38o3vAd9NSM+GFyE0DqNYHzU
M3KgTTrs1ynSDOZ9OFS2OhI5CELfx6qfhmB6z9npyTQm5MOBMG9vp3zoNqGb4i0SqMawBR7JWfbV
uVjS6edoW4K1Dooyz9r3CRUHuOP0Nuiq2VdhFOQ3LeRrAirEYnpS4DgsWxbxI093kX/n59tVMw8r
UJuzUTH/wcjJEbZ95BSCtzkKVi+7Bv14rzQbaikFMHxvzvcBD2YotvQUGiEQMTeCZfJDQHgPnDGe
Egdo63PGlJkqFz9vx+SN59x0F7Cw2nhFeRNm2O4KLaoxpSQRGPOMtvgPMPkK/nUrG8vyKiPk1Yr1
G9GV+3ISuc3EIGP8y7CL2RuQc/yuSsBd3bDuYT/ddqYeEeGYRNkrx5zbJ+SDqNV3nNr6n/vx7cLn
xXhbh4+CH3FMNyRW08dS7vxEhs4H/FzxykWYHbYtO/CReHwRJPg4vaF21WRBtGZEjNcwJPMwRcYO
C/iKpto7mDvZ0tjM0qBCGi4uV2n7PaGtU4fth0YiKy1Oml9e6U2QBVgWkNHUO+QiS2reqlyTvCrE
5VjU+WyV1Z9yTCTZBXAXKJjzbAvVvSS4G29N0Z9YQzVkkpIPXDaP0qEBNUCfPGYcNReCiKMKI4Mz
K9OFFOMiGTVUgtpQOZWcT8J+UvSNPez3gPEaFvumV6lnQvXVX6JZT8WdcXqTbKj9DiNVCHO/dcsJ
MdkM3GwDK3JLt7xVJro3W6eGTcI7LgAB6QIVgc3/aKWjKmbzCys67sHUOkChXl6LpqQN6vUuQxMi
TYlM3X3IkVTW0WqdH7Ht7T6BH8+XZnx0KWi0720LTpsKvqtKGmJfdX3cM3i68NxbgnUVSbnxXrMi
w3bUqdAbSk3VuKSKB8kGTp22JmqlN8+V41CcLAssWls79JeCL0jWmVGvEZwF821KVKo4LoKvahXg
dEwZ2jrGJtuc2+XbY/6Tw83/gJSZhkn9+p/QhIB/RScV3DYpciZj2WT7cIsS74scFWvcbZKmV0qZ
Gd698g4Xeg6YpS4fr9DNx+2INvkeOshlnAYFw7eTtipAQrFDYH45n73+1TozieCSwstZ+yOTZJcX
Niws/ef2UGF2I60zm3O94bs3zTb3U3FqxCRjImw8F8B/HVyBnwh9AJaEikANOg5JuwB1VcB6/vwM
dXtAYqSCT/PIOXqwKXv5+mhk7/j1BokREeP2LcqoJyQqJJZHxW4InH1rq4lO7QRs0qEmWkZTArRo
uCaIjhGUjMNLYSaPEmrhpXlXltNuybJrYtdH2yocB4ItmaRpOmQsACJK9nAxTUgpxsF5NMkKFxmD
Xhb5wdiFDFRGEpSejXQzJvcis4hICfQJn+mtyaq9N7pw3DSIaBMzHbv+Q2c9DoZNrCIh/X9w3MRe
TNaKHv9on5ouSkqujjG/agBJtfIXisRvBP6Lv/o+i8m0XF+E9j6egnHVoYM1D8UhxBRTrji05IkU
p+aK7WcTVcnX7TAxJOUaNZOLeBH04Liboq5oPpvuIHbwFVxm2G4UI4y7uYmnpbp5kHscGnew8Xgp
KM6oSjU5q4uVD5F2nETYCnU47dPZuQB1Hhj/zclt+zQjU0fOLjpq8O4Fck2jpFgXEr8vH5cU4mzp
kLua0/V95FufekuyKrt79XObytu/ZYnCvdJRIsz0umwhM1cqM+GzAMlpfNtGc5NL6Z3wrX3ZFcxO
A5Hj5R/ux1SES1vOHqRrmaJ8bgbfs5egj6qpB58fPet45tJSX/q/wPKNZfzZHACxmVi/cTrDlb/Y
1LPyJrEuPCX1QfTyj0ukGWV7edDZlBHAG7GyWXzcz/aNS2vnQlIjGyI1womSsYYGPeOf+Ij+Ui7i
i/7XtCB83eyzJY5pCednqCsYRh72w1nbMc0qc+v+xIDIHiZ5NrSq0626B4Q+LZG9GiA28fNIhVMz
XDF3EJPmSW2W24RnnT57UfKHJGjgLgCbylreNm5jBa5RJQ3I52McDgIzL8ERd/LgVBxa6+SO0etP
r4JMHAe1u3JX5sTJwtRS2Nq5EMSMA6NhhCvASbHocovsAO7aj9bP1pKBCF1Y15R0aPGo3V48Nj02
AhW7OApEmWUf+tQwThXlu1MK2UGzH5Y8aNygtYPwEZhJKZkLaOhb0YtSBRM4mO8n1e85tSSMyZYL
AD9VvGx55ohdws8wtOyLJP6EW3q3qZOIweSMt5lh0BDLSnKwLTbmxZdOe3+6ntmLvWVrE4+BUBkh
VBHdnr/kKBdkvxTqT5w21TfDZzwuh5f7QYPRXlFpHXeaNsSbTRdttJ+ooRDzRmj86JwURbR+/CzB
xh4tyzRWSpKm+XaftN4IFdBt79lg+meMLuiGBrNlipIlxZ/63uaRsV9E+4MYCDN10y1MwKnBW2c0
mh1aKGkmcBkUdL851z6pb4r3g1GfGSzjoAIkjdEZHT8tD5173KtdqMQ4fSO4Vsm3O8jtwV3LU38I
VGQs21uMa7XA/MhTtFd3sre9eRfBx3fSgoU2r36fKTpvEfq2O917jWQZ8iMOor6xQ6H9UqLEUTNt
AILNf6tcUuYTyA+HCsvHtRwXOMNBg0e1L6FojMN73lZ89DtIcvuXRqa/WbhcteWPm2Y79N2JXcPC
vbDtqIdf71eh5DocDZHcOzwUNX6M087Qfv7gh+4XxVTfKTWm5umcXyb5of78dCHdHj8ZiK01YFjz
qk+J2BBAuT9/FvM9ipr6/jcaxTpFRoM/O74nMk1bdFvjVAsDsGODrcpXMaU8OyOvezBe/GVwyk3A
OqLKONIOXqpMB2Zi6iZHJ1zHp6jHiHH47qmkJD6E77U2y6BuuyvDo8xeGW9XYhc=
`protect end_protected
